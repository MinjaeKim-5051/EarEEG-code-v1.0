`timescale 1 ns/100 ps
// Version: v11.9 SP5 11.9.5.5


module fifo_1b_1b(
       DATA,
       Q,
       WE,
       RE,
       WCLOCK,
       RCLOCK,
       FULL,
       EMPTY,
       RESET,
       RDCNT
    );
input  DATA;
output Q;
input  WE;
input  RE;
input  WCLOCK;
input  RCLOCK;
output FULL;
output EMPTY;
input  RESET;
output [12:0] RDCNT;

    wire RESET_POLA, READ_RESET_P, WRITE_RESET_P, \MEM_RADDR[0] , 
        \RBINNXTSHIFT[0] , \WBINSYNCSHIFT[0] , \MEM_WADDR[0] , 
        \WBINNXTSHIFT[0] , \RBINSYNCSHIFT[0] , \MEM_RADDR[1] , 
        \RBINNXTSHIFT[1] , \WBINSYNCSHIFT[1] , \MEM_WADDR[1] , 
        \WBINNXTSHIFT[1] , \RBINSYNCSHIFT[1] , \MEM_RADDR[2] , 
        \RBINNXTSHIFT[2] , \WBINSYNCSHIFT[2] , \MEM_WADDR[2] , 
        \WBINNXTSHIFT[2] , \RBINSYNCSHIFT[2] , \MEM_RADDR[3] , 
        \RBINNXTSHIFT[3] , \WBINSYNCSHIFT[3] , \MEM_WADDR[3] , 
        \WBINNXTSHIFT[3] , \RBINSYNCSHIFT[3] , \MEM_RADDR[4] , 
        \RBINNXTSHIFT[4] , \WBINSYNCSHIFT[4] , \MEM_WADDR[4] , 
        \WBINNXTSHIFT[4] , \RBINSYNCSHIFT[4] , \MEM_RADDR[5] , 
        \RBINNXTSHIFT[5] , \WBINSYNCSHIFT[5] , \MEM_WADDR[5] , 
        \WBINNXTSHIFT[5] , \RBINSYNCSHIFT[5] , \MEM_RADDR[6] , 
        \RBINNXTSHIFT[6] , \WBINSYNCSHIFT[6] , \MEM_WADDR[6] , 
        \WBINNXTSHIFT[6] , \RBINSYNCSHIFT[6] , \MEM_RADDR[7] , 
        \RBINNXTSHIFT[7] , \WBINSYNCSHIFT[7] , \MEM_WADDR[7] , 
        \WBINNXTSHIFT[7] , \RBINSYNCSHIFT[7] , \MEM_RADDR[8] , 
        \RBINNXTSHIFT[8] , \WBINSYNCSHIFT[8] , \MEM_WADDR[8] , 
        \WBINNXTSHIFT[8] , \RBINSYNCSHIFT[8] , \MEM_RADDR[9] , 
        \RBINNXTSHIFT[9] , \WBINSYNCSHIFT[9] , \MEM_WADDR[9] , 
        \WBINNXTSHIFT[9] , \RBINSYNCSHIFT[9] , \MEM_RADDR[10] , 
        \RBINNXTSHIFT[10] , \WBINSYNCSHIFT[10] , \MEM_WADDR[10] , 
        \WBINNXTSHIFT[10] , \RBINSYNCSHIFT[10] , \MEM_RADDR[11] , 
        \RBINNXTSHIFT[11] , \WBINSYNCSHIFT[11] , \MEM_WADDR[11] , 
        \WBINNXTSHIFT[11] , \RBINSYNCSHIFT[11] , \MEM_RADDR[12] , 
        \RBINNXTSHIFT[12] , READDOMAIN_WMSB, \MEM_WADDR[12] , 
        \WBINNXTSHIFT[12] , \RBINSYNCSHIFT[12] , FULLINT, MEMORYWE, 
        MEMWENEG, \WGRY[0] , \WGRY[1] , \WGRY[2] , \WGRY[3] , 
        \WGRY[4] , \WGRY[5] , \WGRY[6] , \WGRY[7] , \WGRY[8] , 
        \WGRY[9] , \WGRY[10] , \WGRY[11] , \WGRY[12] , \RGRYSYNC[0] , 
        \RGRYSYNC[1] , \RGRYSYNC[2] , \RGRYSYNC[3] , \RGRYSYNC[4] , 
        \RGRYSYNC[5] , \RGRYSYNC[6] , \RGRYSYNC[7] , \RGRYSYNC[8] , 
        \RGRYSYNC[9] , \RGRYSYNC[10] , \RGRYSYNC[11] , \RGRYSYNC[12] , 
        EMPTYINT, MEMORYRE, MEMRENEG, \RDIFF[0] , \RDIFF[1] , 
        \RDIFF[2] , \RDIFF[3] , \RDIFF[4] , \RDIFF[5] , \RDIFF[6] , 
        \RDIFF[7] , \RDIFF[8] , \RDIFF[9] , \RDIFF[10] , \RDIFF[11] , 
        \RDIFF[12] , DVLDI, DVLDX, \RGRY[0] , \RGRY[1] , \RGRY[2] , 
        \RGRY[3] , \RGRY[4] , \RGRY[5] , \RGRY[6] , \RGRY[7] , 
        \RGRY[8] , \RGRY[9] , \RGRY[10] , \RGRY[11] , \RGRY[12] , 
        \WGRYSYNC[0] , \WGRYSYNC[1] , \WGRYSYNC[2] , \WGRYSYNC[3] , 
        \WGRYSYNC[4] , \WGRYSYNC[5] , \WGRYSYNC[6] , \WGRYSYNC[7] , 
        \WGRYSYNC[8] , \WGRYSYNC[9] , \WGRYSYNC[10] , \WGRYSYNC[11] , 
        \WGRYSYNC[12] , QXI, NOR2A_0_Y, INV_0_Y, INV_9_Y, INV_2_Y, 
        INV_12_Y, INV_10_Y, INV_5_Y, INV_7_Y, INV_1_Y, INV_3_Y, 
        INV_11_Y, INV_8_Y, INV_6_Y, INV_4_Y, AND2_37_Y, AND2_22_Y, 
        AND2_67_Y, AND2_55_Y, AND2_92_Y, AND2_51_Y, AND2_53_Y, 
        AND2_90_Y, AND2_74_Y, AND2_50_Y, AND2_60_Y, AND2_59_Y, 
        AND2_35_Y, AND2_48_Y, XOR2_10_Y, XOR2_11_Y, XOR2_0_Y, 
        XOR2_49_Y, XOR2_19_Y, XOR2_44_Y, XOR2_41_Y, XOR2_94_Y, 
        XOR2_14_Y, XOR2_91_Y, XOR2_26_Y, XOR2_82_Y, AND2_12_Y, 
        AO1_10_Y, AND2_21_Y, AO1_23_Y, AND2_8_Y, AO1_13_Y, AND2_30_Y, 
        AO1_44_Y, AND2_88_Y, AO1_11_Y, AND2_42_Y, AND2_96_Y, AO1_19_Y, 
        AND2_80_Y, AO1_43_Y, AND2_63_Y, AND2_75_Y, AO1_38_Y, AND2_6_Y, 
        AND2_15_Y, AND2_2_Y, AND2_23_Y, AND2_77_Y, AND2_32_Y, 
        AND2_89_Y, AND2_72_Y, OR3_0_Y, AO1_4_Y, AO1_53_Y, AO1_2_Y, 
        AO1_52_Y, AO1_28_Y, AO1_14_Y, AO1_5_Y, AO1_51_Y, AO1_41_Y, 
        AO1_3_Y, XOR2_89_Y, XOR2_32_Y, XOR2_51_Y, XOR2_64_Y, XOR2_29_Y, 
        XOR2_93_Y, XOR2_38_Y, XOR2_60_Y, XOR2_72_Y, XOR2_48_Y, 
        XOR2_12_Y, XOR2_61_Y, DFN1C0_13_Q, DFN1C0_10_Q, DFN1C0_11_Q, 
        DFN1C0_26_Q, DFN1C0_5_Q, DFN1C0_24_Q, DFN1C0_20_Q, DFN1C0_8_Q, 
        DFN1C0_23_Q, DFN1C0_22_Q, DFN1C0_2_Q, DFN1C0_12_Q, DFN1C0_17_Q, 
        XNOR3_1_Y, XNOR3_39_Y, XOR3_2_Y, XNOR3_47_Y, XNOR3_46_Y, 
        XNOR3_0_Y, XOR3_5_Y, XNOR3_24_Y, XNOR3_51_Y, XOR3_1_Y, 
        XNOR3_42_Y, XNOR3_45_Y, XNOR3_10_Y, XNOR3_3_Y, XNOR3_44_Y, 
        XOR3_7_Y, XNOR3_49_Y, XNOR3_7_Y, XNOR3_19_Y, XNOR3_2_Y, 
        XNOR3_37_Y, XNOR3_36_Y, XNOR3_41_Y, XNOR3_9_Y, XNOR3_30_Y, 
        XNOR3_23_Y, XNOR3_43_Y, XNOR3_12_Y, XNOR3_6_Y, XNOR3_5_Y, 
        XOR2_18_Y, XOR2_28_Y, XOR2_57_Y, XOR2_58_Y, XOR2_84_Y, 
        XOR2_92_Y, XOR2_75_Y, XOR2_24_Y, XOR2_74_Y, XOR2_43_Y, 
        XOR2_87_Y, XOR2_6_Y, XOR2_45_Y, AND2_49_Y, AND2_20_Y, 
        AND2_68_Y, AND2_5_Y, AND2_19_Y, AND2_1_Y, AND2_43_Y, AND2_34_Y, 
        AND2_46_Y, AND2_38_Y, AND2_45_Y, AND2_84_Y, XOR2_76_Y, 
        XOR2_7_Y, XOR2_13_Y, XOR2_4_Y, XOR2_15_Y, XOR2_31_Y, XOR2_71_Y, 
        XOR2_5_Y, XOR2_20_Y, XOR2_85_Y, XOR2_68_Y, XOR2_8_Y, XOR2_95_Y, 
        AND2_24_Y, AO1_45_Y, AND2_79_Y, AO1_16_Y, AND2_27_Y, AO1_55_Y, 
        AND2_44_Y, AO1_47_Y, AND2_70_Y, AO1_25_Y, AND2_61_Y, AND2_87_Y, 
        AO1_48_Y, AND2_4_Y, AO1_0_Y, AND2_83_Y, AND2_0_Y, AND2_94_Y, 
        AND2_52_Y, AND2_95_Y, AND2_16_Y, AND2_47_Y, AND2_40_Y, 
        AND2_56_Y, AND2_93_Y, AO1_46_Y, AND2_69_Y, AND2_91_Y, AO1_24_Y, 
        AO1_35_Y, AO1_12_Y, AO1_20_Y, AO1_6_Y, AO1_32_Y, AO1_29_Y, 
        AO1_15_Y, AO1_26_Y, AO1_54_Y, AO1_49_Y, XOR2_50_Y, XOR2_46_Y, 
        XOR2_69_Y, XOR2_96_Y, XOR2_27_Y, XOR2_88_Y, XOR2_83_Y, 
        XOR2_97_Y, XOR2_9_Y, XOR2_39_Y, XOR2_100_Y, XOR2_98_Y, 
        NAND2_1_Y, XOR2_42_Y, XOR2_35_Y, XOR2_23_Y, XOR2_73_Y, 
        XOR2_63_Y, XOR2_37_Y, XOR2_52_Y, XOR2_59_Y, XOR2_62_Y, 
        XOR2_21_Y, XOR2_54_Y, XOR2_3_Y, XOR2_70_Y, AND2_66_Y, 
        AND2_13_Y, AND2_9_Y, AND2_71_Y, AND2_14_Y, AND2_78_Y, 
        AND2_18_Y, AND2_85_Y, AND2_73_Y, AND2_3_Y, AND2_7_Y, AND2_33_Y, 
        XOR2_47_Y, XOR2_40_Y, XOR2_22_Y, XOR2_86_Y, XOR2_81_Y, 
        XOR2_77_Y, XOR2_1_Y, XOR2_65_Y, XOR2_25_Y, XOR2_56_Y, 
        XOR2_79_Y, XOR2_30_Y, XOR2_34_Y, AND2_82_Y, AO1_31_Y, 
        AND2_81_Y, AO1_7_Y, AND2_86_Y, AO1_8_Y, AND2_65_Y, AO1_27_Y, 
        AND2_11_Y, AO1_50_Y, AND2_17_Y, AND2_41_Y, AO1_34_Y, AND2_36_Y, 
        AO1_40_Y, AND2_64_Y, AND2_58_Y, AND2_29_Y, AND2_28_Y, 
        AND2_31_Y, AND2_10_Y, AND2_54_Y, AND2_62_Y, AND2_76_Y, 
        AND2_26_Y, AO1_33_Y, AND2_57_Y, AND2_39_Y, AO1_1_Y, AO1_37_Y, 
        AO1_36_Y, AO1_30_Y, AO1_17_Y, AO1_18_Y, AO1_9_Y, AO1_39_Y, 
        AO1_21_Y, AO1_42_Y, AO1_22_Y, XOR2_66_Y, XOR2_16_Y, XOR2_90_Y, 
        XOR2_99_Y, XOR2_53_Y, XOR2_78_Y, XOR2_33_Y, XOR2_2_Y, 
        XOR2_80_Y, XOR2_36_Y, XOR2_67_Y, XOR2_17_Y, XNOR3_27_Y, 
        XNOR3_8_Y, XOR3_0_Y, XNOR3_18_Y, XNOR3_22_Y, XNOR3_26_Y, 
        XOR3_3_Y, XNOR3_50_Y, XNOR3_25_Y, XOR3_6_Y, XNOR3_14_Y, 
        XNOR3_21_Y, XNOR3_33_Y, XNOR3_29_Y, XNOR3_16_Y, XOR3_4_Y, 
        XNOR3_20_Y, XNOR3_31_Y, XNOR3_38_Y, XNOR3_28_Y, XNOR3_17_Y, 
        XNOR3_40_Y, XNOR3_13_Y, XNOR3_32_Y, XNOR3_4_Y, XNOR3_48_Y, 
        XNOR3_15_Y, XNOR3_34_Y, XNOR3_35_Y, XNOR3_11_Y, DFN1C0_27_Q, 
        DFN1C0_0_Q, DFN1C0_6_Q, DFN1C0_18_Q, DFN1C0_4_Q, DFN1C0_14_Q, 
        DFN1C0_21_Q, DFN1C0_16_Q, DFN1C0_25_Q, DFN1C0_1_Q, DFN1C0_7_Q, 
        DFN1C0_9_Q, DFN1C0_19_Q, RAM4K9_QXI_DOUTA0, AND3_0_Y, 
        XNOR2_22_Y, XNOR2_12_Y, XNOR2_7_Y, XNOR2_13_Y, XNOR2_14_Y, 
        XNOR2_24_Y, XNOR2_10_Y, XNOR2_18_Y, XNOR2_20_Y, XNOR2_16_Y, 
        XNOR2_9_Y, XNOR2_23_Y, XNOR2_4_Y, AND3_7_Y, AND3_8_Y, 
        AND2_25_Y, AND3_9_Y, AND3_6_Y, DFN1C0_15_Q, AND2A_0_Y, 
        DFN1C0_3_Q, AND3_1_Y, XOR2_55_Y, XNOR2_1_Y, XNOR2_17_Y, 
        XNOR2_21_Y, XNOR2_19_Y, XNOR2_0_Y, XNOR2_5_Y, XNOR2_15_Y, 
        XNOR2_8_Y, XNOR2_2_Y, XNOR2_3_Y, XNOR2_6_Y, XNOR2_11_Y, 
        AND3_5_Y, AND3_2_Y, AND2_97_Y, AND3_4_Y, AND3_3_Y, NAND2_0_Y, 
        VCC, GND;
    wire GND_power_net1;
    wire VCC_power_net1;
    assign GND = GND_power_net1;
    assign VCC = VCC_power_net1;
    
    DFN1C0 \DFN1C0_RDCNT[2]  (.D(\RDIFF[2] ), .CLK(RCLOCK), .CLR(
        READ_RESET_P), .Q(RDCNT[2]));
    XNOR3 XNOR3_14 (.A(\WGRYSYNC[9] ), .B(\WGRYSYNC[8] ), .C(
        \WGRYSYNC[7] ), .Y(XNOR3_14_Y));
    INV INV_0 (.A(\RBINNXTSHIFT[1] ), .Y(INV_0_Y));
    AO1 AO1_52 (.A(XOR2_19_Y), .B(AO1_2_Y), .C(AND2_53_Y), .Y(AO1_52_Y)
        );
    XNOR3 XNOR3_5 (.A(\RGRYSYNC[0] ), .B(XNOR3_6_Y), .C(XNOR3_23_Y), 
        .Y(XNOR3_5_Y));
    DFN1C0 \DFN1C0_RGRYSYNC[4]  (.D(DFN1C0_4_Q), .CLK(WCLOCK), .CLR(
        WRITE_RESET_P), .Q(\RGRYSYNC[4] ));
    XNOR3 XNOR3_45 (.A(\RGRYSYNC[12] ), .B(\RGRYSYNC[11] ), .C(
        \RGRYSYNC[10] ), .Y(XNOR3_45_Y));
    AND2 AND2_2 (.A(AND2_75_Y), .B(AND2_88_Y), .Y(AND2_2_Y));
    AND3 AND3_6 (.A(XNOR2_14_Y), .B(XNOR2_24_Y), .C(XNOR2_10_Y), .Y(
        AND3_6_Y));
    XOR3 \XOR3_WBINSYNCSHIFT[10]  (.A(\WGRYSYNC[12] ), .B(
        \WGRYSYNC[11] ), .C(\WGRYSYNC[10] ), .Y(\WBINSYNCSHIFT[10] ));
    AND2 AND2_20 (.A(\MEM_RADDR[2] ), .B(GND), .Y(AND2_20_Y));
    XOR2 XOR2_82 (.A(READDOMAIN_WMSB), .B(INV_6_Y), .Y(XOR2_82_Y));
    XNOR2 XNOR2_13 (.A(\RBINNXTSHIFT[2] ), .B(\WBINSYNCSHIFT[2] ), .Y(
        XNOR2_13_Y));
    DFN1C0 \DFN1C0_RDCNT[5]  (.D(\RDIFF[5] ), .CLK(RCLOCK), .CLR(
        READ_RESET_P), .Q(RDCNT[5]));
    AO1 AO1_11 (.A(XOR2_82_Y), .B(AND2_35_Y), .C(AND2_48_Y), .Y(
        AO1_11_Y));
    AND2 AND2_11 (.A(XOR2_25_Y), .B(XOR2_56_Y), .Y(AND2_11_Y));
    XOR2 \XOR2_WBINNXTSHIFT[2]  (.A(XOR2_16_Y), .B(AO1_1_Y), .Y(
        \WBINNXTSHIFT[2] ));
    XNOR3 XNOR3_34 (.A(\WGRYSYNC[3] ), .B(\WGRYSYNC[2] ), .C(
        \WGRYSYNC[1] ), .Y(XNOR3_34_Y));
    XNOR3 XNOR3_25 (.A(\WGRYSYNC[9] ), .B(\WGRYSYNC[8] ), .C(
        \WGRYSYNC[7] ), .Y(XNOR3_25_Y));
    AND2 AND2_22 (.A(\WBINSYNCSHIFT[1] ), .B(INV_4_Y), .Y(AND2_22_Y));
    DFN1C0 \DFN1C0_RGRY[9]  (.D(XOR2_43_Y), .CLK(RCLOCK), .CLR(
        READ_RESET_P), .Q(\RGRY[9] ));
    DFN1C0 DFN1C0_FULL (.D(FULLINT), .CLK(WCLOCK), .CLR(WRITE_RESET_P), 
        .Q(FULL));
    XNOR2 XNOR2_9 (.A(\RBINNXTSHIFT[9] ), .B(\WBINSYNCSHIFT[9] ), .Y(
        XNOR2_9_Y));
    XOR3 \XOR3_RBINSYNCSHIFT[10]  (.A(\RGRYSYNC[12] ), .B(
        \RGRYSYNC[11] ), .C(\RGRYSYNC[10] ), .Y(\RBINSYNCSHIFT[10] ));
    AND2 AND2_71 (.A(\MEM_WADDR[4] ), .B(GND), .Y(AND2_71_Y));
    DFN1C0 DFN1C0_17 (.D(\WGRY[12] ), .CLK(RCLOCK), .CLR(READ_RESET_P), 
        .Q(DFN1C0_17_Q));
    XOR2 XOR2_19 (.A(\WBINSYNCSHIFT[5] ), .B(INV_10_Y), .Y(XOR2_19_Y));
    AND2 AND2_44 (.A(XOR2_71_Y), .B(XOR2_5_Y), .Y(AND2_44_Y));
    AO1 AO1_31 (.A(XOR2_86_Y), .B(AND2_13_Y), .C(AND2_9_Y), .Y(
        AO1_31_Y));
    DFN1C0 \DFN1C0_RDCNT[12]  (.D(\RDIFF[12] ), .CLK(RCLOCK), .CLR(
        READ_RESET_P), .Q(RDCNT[12]));
    XOR2 XOR2_1 (.A(\MEM_WADDR[6] ), .B(GND), .Y(XOR2_1_Y));
    XOR2 XOR2_23 (.A(\WBINNXTSHIFT[2] ), .B(\WBINNXTSHIFT[3] ), .Y(
        XOR2_23_Y));
    XOR2 XOR2_100 (.A(\MEM_RADDR[11] ), .B(GND), .Y(XOR2_100_Y));
    XNOR3 XNOR3_13 (.A(\WGRYSYNC[9] ), .B(\WGRYSYNC[8] ), .C(
        \WGRYSYNC[7] ), .Y(XNOR3_13_Y));
    DFN1C0 \DFN1C0_RGRYSYNC[3]  (.D(DFN1C0_18_Q), .CLK(WCLOCK), .CLR(
        WRITE_RESET_P), .Q(\RGRYSYNC[3] ));
    XOR2 \XOR2_RDIFF[10]  (.A(XOR2_48_Y), .B(AO1_51_Y), .Y(\RDIFF[10] )
        );
    INV INV_1 (.A(\RBINNXTSHIFT[8] ), .Y(INV_1_Y));
    XOR2 XOR2_47 (.A(\MEM_WADDR[0] ), .B(MEMORYWE), .Y(XOR2_47_Y));
    XOR2 XOR2_38 (.A(\WBINSYNCSHIFT[7] ), .B(INV_7_Y), .Y(XOR2_38_Y));
    BUFF BUFF_READDOMAIN_WMSB (.A(\WGRYSYNC[12] ), .Y(READDOMAIN_WMSB));
    XOR2 \XOR2_RBINNXTSHIFT[0]  (.A(\MEM_RADDR[0] ), .B(MEMORYRE), .Y(
        \RBINNXTSHIFT[0] ));
    AO1 AO1_7 (.A(XOR2_77_Y), .B(AND2_71_Y), .C(AND2_14_Y), .Y(AO1_7_Y)
        );
    DFN1C0 DFN1C0_9 (.D(\RGRY[11] ), .CLK(WCLOCK), .CLR(WRITE_RESET_P), 
        .Q(DFN1C0_9_Q));
    DFN1C0 \DFN1C0_WGRY[6]  (.D(XOR2_52_Y), .CLK(WCLOCK), .CLR(
        WRITE_RESET_P), .Q(\WGRY[6] ));
    AND2 AND2_18 (.A(\MEM_WADDR[7] ), .B(GND), .Y(AND2_18_Y));
    AND2 AND2_15 (.A(AND2_96_Y), .B(AND2_8_Y), .Y(AND2_15_Y));
    AND2 AND2_84 (.A(\MEM_RADDR[12] ), .B(GND), .Y(AND2_84_Y));
    XNOR3 XNOR3_33 (.A(\WGRYSYNC[6] ), .B(\WGRYSYNC[5] ), .C(
        XNOR3_21_Y), .Y(XNOR3_33_Y));
    DFN1C0 DFN1C0_WRITE_RESET_P (.D(DFN1C0_15_Q), .CLK(WCLOCK), .CLR(
        RESET_POLA), .Q(WRITE_RESET_P));
    INV INV_7 (.A(\RBINNXTSHIFT[7] ), .Y(INV_7_Y));
    AO1 AO1_25 (.A(XOR2_8_Y), .B(AND2_38_Y), .C(AND2_45_Y), .Y(
        AO1_25_Y));
    DFN1C0 DFN1C0_26 (.D(\WGRY[3] ), .CLK(RCLOCK), .CLR(READ_RESET_P), 
        .Q(DFN1C0_26_Q));
    AND2 AND2_78 (.A(\MEM_WADDR[6] ), .B(GND), .Y(AND2_78_Y));
    AND2 AND2_75 (.A(AND2_96_Y), .B(AND2_80_Y), .Y(AND2_75_Y));
    XOR2 \XOR2_RDIFF[3]  (.A(XOR2_51_Y), .B(AO1_4_Y), .Y(\RDIFF[3] ));
    XOR2 XOR2_45 (.A(\RBINNXTSHIFT[12] ), .B(GND), .Y(XOR2_45_Y));
    DFN1C0 \DFN1C0_RGRYSYNC[7]  (.D(DFN1C0_16_Q), .CLK(WCLOCK), .CLR(
        WRITE_RESET_P), .Q(\RGRYSYNC[7] ));
    XOR2 \XOR2_RBINNXTSHIFT[9]  (.A(XOR2_9_Y), .B(AO1_15_Y), .Y(
        \RBINNXTSHIFT[9] ));
    DFN1C0 DFN1C0_11 (.D(\WGRY[2] ), .CLK(RCLOCK), .CLR(READ_RESET_P), 
        .Q(DFN1C0_11_Q));
    DFN1C0 DFN1C0_0 (.D(\RGRY[1] ), .CLK(WCLOCK), .CLR(WRITE_RESET_P), 
        .Q(DFN1C0_0_Q));
    BUFF \BUFF_RBINSYNCSHIFT[12]  (.A(\RGRYSYNC[12] ), .Y(
        \RBINSYNCSHIFT[12] ));
    AND2 AND2_1 (.A(\MEM_RADDR[6] ), .B(GND), .Y(AND2_1_Y));
    DFN1C0 \DFN1C0_MEM_WADDR[0]  (.D(\WBINNXTSHIFT[0] ), .CLK(WCLOCK), 
        .CLR(WRITE_RESET_P), .Q(\MEM_WADDR[0] ));
    XNOR2 XNOR2_21 (.A(\RBINSYNCSHIFT[2] ), .B(\WBINNXTSHIFT[2] ), .Y(
        XNOR2_21_Y));
    DFN1C0 \DFN1C0_MEM_WADDR[3]  (.D(\WBINNXTSHIFT[3] ), .CLK(WCLOCK), 
        .CLR(WRITE_RESET_P), .Q(\MEM_WADDR[3] ));
    AND2 AND2_49 (.A(\MEM_RADDR[1] ), .B(GND), .Y(AND2_49_Y));
    DFN1C0 \DFN1C0_MEM_RADDR[1]  (.D(\RBINNXTSHIFT[1] ), .CLK(RCLOCK), 
        .CLR(READ_RESET_P), .Q(\MEM_RADDR[1] ));
    AO1 AO1_8 (.A(XOR2_65_Y), .B(AND2_78_Y), .C(AND2_18_Y), .Y(AO1_8_Y)
        );
    DFN1C0 DFN1C0_20 (.D(\WGRY[6] ), .CLK(RCLOCK), .CLR(READ_RESET_P), 
        .Q(DFN1C0_20_Q));
    AND2 AND2_10 (.A(AND2_82_Y), .B(XOR2_22_Y), .Y(AND2_10_Y));
    XOR2 XOR2_92 (.A(\RBINNXTSHIFT[5] ), .B(\RBINNXTSHIFT[6] ), .Y(
        XOR2_92_Y));
    DFN1C0 \DFN1C0_RGRYSYNC[6]  (.D(DFN1C0_21_Q), .CLK(WCLOCK), .CLR(
        WRITE_RESET_P), .Q(\RGRYSYNC[6] ));
    AND2 AND2_7 (.A(\MEM_WADDR[11] ), .B(GND), .Y(AND2_7_Y));
    XOR2 XOR2_20 (.A(\MEM_RADDR[8] ), .B(GND), .Y(XOR2_20_Y));
    XOR2 XOR2_63 (.A(\WBINNXTSHIFT[4] ), .B(\WBINNXTSHIFT[5] ), .Y(
        XOR2_63_Y));
    XOR2 XOR2_87 (.A(\RBINNXTSHIFT[10] ), .B(\RBINNXTSHIFT[11] ), .Y(
        XOR2_87_Y));
    AND2 AND2_70 (.A(XOR2_20_Y), .B(XOR2_85_Y), .Y(AND2_70_Y));
    AND2 AND2_12 (.A(XOR2_10_Y), .B(XOR2_11_Y), .Y(AND2_12_Y));
    DFN1C0 \DFN1C0_WGRY[5]  (.D(XOR2_37_Y), .CLK(WCLOCK), .CLR(
        WRITE_RESET_P), .Q(\WGRY[5] ));
    AO1 AO1_42 (.A(XOR2_79_Y), .B(AO1_21_Y), .C(AND2_3_Y), .Y(AO1_42_Y)
        );
    XOR2 XOR2_52 (.A(\WBINNXTSHIFT[6] ), .B(\WBINNXTSHIFT[7] ), .Y(
        XOR2_52_Y));
    XNOR3 XNOR3_40 (.A(XNOR3_17_Y), .B(XNOR3_31_Y), .C(XNOR3_38_Y), .Y(
        XNOR3_40_Y));
    XOR2 \XOR2_WBINNXTSHIFT[0]  (.A(\MEM_WADDR[0] ), .B(MEMORYWE), .Y(
        \WBINNXTSHIFT[0] ));
    AO1 AO1_50 (.A(XOR2_30_Y), .B(AND2_3_Y), .C(AND2_7_Y), .Y(AO1_50_Y)
        );
    AND2 AND2_72 (.A(AND2_2_Y), .B(XOR2_26_Y), .Y(AND2_72_Y));
    DFN1C0 \DFN1C0_MEM_WADDR[4]  (.D(\WBINNXTSHIFT[4] ), .CLK(WCLOCK), 
        .CLR(WRITE_RESET_P), .Q(\MEM_WADDR[4] ));
    AND2 AND2_61 (.A(XOR2_68_Y), .B(XOR2_8_Y), .Y(AND2_61_Y));
    AO1 AO1_15 (.A(XOR2_20_Y), .B(AO1_29_Y), .C(AND2_34_Y), .Y(
        AO1_15_Y));
    DFN1C0 \DFN1C0_WGRY[7]  (.D(XOR2_59_Y), .CLK(WCLOCK), .CLR(
        WRITE_RESET_P), .Q(\WGRY[7] ));
    DFN1C0 \DFN1C0_MEM_WADDR[12]  (.D(\WBINNXTSHIFT[12] ), .CLK(WCLOCK)
        , .CLR(WRITE_RESET_P), .Q(\MEM_WADDR[12] ));
    DFN1C0 DFN1C0_READ_RESET_P (.D(DFN1C0_3_Q), .CLK(RCLOCK), .CLR(
        RESET_POLA), .Q(READ_RESET_P));
    XNOR3 \XNOR3_WBINSYNCSHIFT[2]  (.A(XNOR3_29_Y), .B(XNOR3_16_Y), .C(
        XNOR3_20_Y), .Y(\WBINSYNCSHIFT[2] ));
    AND2 AND2_EMPTYINT (.A(AND3_0_Y), .B(XNOR2_22_Y), .Y(EMPTYINT));
    XOR2 XOR2_85 (.A(\MEM_RADDR[9] ), .B(GND), .Y(XOR2_85_Y));
    XNOR2 \XNOR2_RBINSYNCSHIFT[5]  (.A(XNOR3_42_Y), .B(XNOR3_10_Y), .Y(
        \RBINSYNCSHIFT[5] ));
    AND2 AND2_89 (.A(AND2_75_Y), .B(XOR2_14_Y), .Y(AND2_89_Y));
    XOR2 XOR2_24 (.A(\RBINNXTSHIFT[7] ), .B(\RBINNXTSHIFT[8] ), .Y(
        XOR2_24_Y));
    AND2 AND2_57 (.A(AND2_29_Y), .B(XOR2_34_Y), .Y(AND2_57_Y));
    XNOR3 XNOR3_20 (.A(\WGRYSYNC[3] ), .B(\WGRYSYNC[2] ), .C(XOR3_4_Y), 
        .Y(XNOR3_20_Y));
    XOR2 XOR2_21 (.A(\WBINNXTSHIFT[9] ), .B(\WBINNXTSHIFT[10] ), .Y(
        XOR2_21_Y));
    AO1 AO1_35 (.A(XOR2_13_Y), .B(AO1_24_Y), .C(AND2_20_Y), .Y(
        AO1_35_Y));
    XOR2 \XOR2_WBINNXTSHIFT[9]  (.A(XOR2_80_Y), .B(AO1_39_Y), .Y(
        \WBINNXTSHIFT[9] ));
    DFN1C0 \DFN1C0_WGRYSYNC[11]  (.D(DFN1C0_12_Q), .CLK(RCLOCK), .CLR(
        READ_RESET_P), .Q(\WGRYSYNC[11] ));
    XNOR2 \XNOR2_RBINSYNCSHIFT[9]  (.A(\RGRYSYNC[9] ), .B(XNOR3_46_Y), 
        .Y(\RBINSYNCSHIFT[9] ));
    DFN1C0 \DFN1C0_WGRYSYNC[12]  (.D(DFN1C0_17_Q), .CLK(RCLOCK), .CLR(
        READ_RESET_P), .Q(\WGRYSYNC[12] ));
    INV INV_11 (.A(\RBINNXTSHIFT[10] ), .Y(INV_11_Y));
    AND2 AND2_46 (.A(\MEM_RADDR[9] ), .B(GND), .Y(AND2_46_Y));
    AO1 AO1_53 (.A(XOR2_0_Y), .B(AO1_4_Y), .C(AND2_92_Y), .Y(AO1_53_Y));
    XNOR3 XNOR3_9 (.A(\RGRYSYNC[6] ), .B(\RGRYSYNC[5] ), .C(
        \RGRYSYNC[4] ), .Y(XNOR3_9_Y));
    XNOR3 XNOR3_8 (.A(\WGRYSYNC[6] ), .B(\WGRYSYNC[5] ), .C(
        \WGRYSYNC[4] ), .Y(XNOR3_8_Y));
    XOR2 \XOR2_RBINNXTSHIFT[8]  (.A(XOR2_97_Y), .B(AO1_29_Y), .Y(
        \RBINNXTSHIFT[8] ));
    XNOR2 \XNOR2_RBINSYNCSHIFT[1]  (.A(XNOR3_2_Y), .B(XNOR3_36_Y), .Y(
        \RBINSYNCSHIFT[1] ));
    XNOR3 XNOR3_50 (.A(\WGRYSYNC[12] ), .B(\WGRYSYNC[11] ), .C(
        \WGRYSYNC[10] ), .Y(XNOR3_50_Y));
    XOR2 XOR2_16 (.A(\MEM_WADDR[2] ), .B(GND), .Y(XOR2_16_Y));
    DFN1C0 DFN1C0_4 (.D(\RGRY[4] ), .CLK(WCLOCK), .CLR(WRITE_RESET_P), 
        .Q(DFN1C0_4_Q));
    XOR2 XOR2_60 (.A(\WBINSYNCSHIFT[8] ), .B(INV_1_Y), .Y(XOR2_60_Y));
    DFN1C0 DFN1C0_14 (.D(\RGRY[5] ), .CLK(WCLOCK), .CLR(WRITE_RESET_P), 
        .Q(DFN1C0_14_Q));
    AND2 AND2_68 (.A(\MEM_RADDR[3] ), .B(GND), .Y(AND2_68_Y));
    AND2 AND2_65 (.A(XOR2_1_Y), .B(XOR2_65_Y), .Y(AND2_65_Y));
    AND2 AND2_43 (.A(\MEM_RADDR[7] ), .B(GND), .Y(AND2_43_Y));
    AO1 AO1_24 (.A(XOR2_7_Y), .B(AND2_91_Y), .C(AND2_49_Y), .Y(
        AO1_24_Y));
    XNOR3 \XNOR3_WBINSYNCSHIFT[8]  (.A(\WGRYSYNC[9] ), .B(
        \WGRYSYNC[8] ), .C(XNOR3_50_Y), .Y(\WBINSYNCSHIFT[8] ));
    AND3 AND3_3 (.A(XNOR2_19_Y), .B(XNOR2_0_Y), .C(XNOR2_5_Y), .Y(
        AND3_3_Y));
    INV INV_5 (.A(\RBINNXTSHIFT[6] ), .Y(INV_5_Y));
    AND2 AND2_86 (.A(XOR2_81_Y), .B(XOR2_77_Y), .Y(AND2_86_Y));
    INV MEMWEBUBBLE (.A(MEMORYWE), .Y(MEMWENEG));
    AND2 AND2_6 (.A(AND2_75_Y), .B(AND2_63_Y), .Y(AND2_6_Y));
    XOR2 XOR2_97 (.A(\MEM_RADDR[8] ), .B(GND), .Y(XOR2_97_Y));
    XOR2 XOR2_64 (.A(\WBINSYNCSHIFT[4] ), .B(INV_12_Y), .Y(XOR2_64_Y));
    AND3 AND3_0 (.A(XNOR2_9_Y), .B(AND3_8_Y), .C(AND2_25_Y), .Y(
        AND3_0_Y));
    DFN1C0 \DFN1C0_MEM_RADDR[2]  (.D(\RBINNXTSHIFT[2] ), .CLK(RCLOCK), 
        .CLR(READ_RESET_P), .Q(\MEM_RADDR[2] ));
    AND2 AND2_60 (.A(\WBINSYNCSHIFT[9] ), .B(INV_3_Y), .Y(AND2_60_Y));
    DFN1C0 \DFN1C0_RGRYSYNC[11]  (.D(DFN1C0_9_Q), .CLK(WCLOCK), .CLR(
        WRITE_RESET_P), .Q(\RGRYSYNC[11] ));
    XOR2 XOR2_61 (.A(READDOMAIN_WMSB), .B(INV_6_Y), .Y(XOR2_61_Y));
    AND2 AND2_83 (.A(AND2_70_Y), .B(AND2_61_Y), .Y(AND2_83_Y));
    XOR2 XOR2_57 (.A(\RBINNXTSHIFT[2] ), .B(\RBINNXTSHIFT[3] ), .Y(
        XOR2_57_Y));
    DFN1C0 \DFN1C0_RGRY[2]  (.D(XOR2_57_Y), .CLK(RCLOCK), .CLR(
        READ_RESET_P), .Q(\RGRY[2] ));
    AND2 AND2_62 (.A(AND2_28_Y), .B(XOR2_1_Y), .Y(AND2_62_Y));
    INV INV_3 (.A(\RBINNXTSHIFT[9] ), .Y(INV_3_Y));
    XOR2 XOR2_33 (.A(\MEM_WADDR[7] ), .B(GND), .Y(XOR2_33_Y));
    AND2 AND2_97 (.A(XNOR2_6_Y), .B(XNOR2_11_Y), .Y(AND2_97_Y));
    XNOR2 XNOR2_2 (.A(\RBINSYNCSHIFT[8] ), .B(\WBINNXTSHIFT[8] ), .Y(
        XNOR2_2_Y));
    XNOR2 XNOR2_19 (.A(\RBINSYNCSHIFT[3] ), .B(\WBINNXTSHIFT[3] ), .Y(
        XNOR2_19_Y));
    XOR2 XOR2_49 (.A(\WBINSYNCSHIFT[4] ), .B(INV_12_Y), .Y(XOR2_49_Y));
    XOR2 \XOR2_WBINNXTSHIFT[8]  (.A(XOR2_2_Y), .B(AO1_9_Y), .Y(
        \WBINNXTSHIFT[8] ));
    XOR2 XOR2_95 (.A(\MEM_RADDR[12] ), .B(GND), .Y(XOR2_95_Y));
    AO1 AO1_14 (.A(XOR2_41_Y), .B(AO1_28_Y), .C(AND2_74_Y), .Y(
        AO1_14_Y));
    XOR2 XOR2_4 (.A(\MEM_RADDR[3] ), .B(GND), .Y(XOR2_4_Y));
    XNOR2 \XNOR2_WBINSYNCSHIFT[3]  (.A(XNOR3_8_Y), .B(XNOR3_18_Y), .Y(
        \WBINSYNCSHIFT[3] ));
    AND3 AND3_1 (.A(XNOR2_3_Y), .B(AND3_2_Y), .C(AND2_97_Y), .Y(
        AND3_1_Y));
    XOR2 XOR2_55 (.A(\RBINSYNCSHIFT[12] ), .B(\WBINNXTSHIFT[12] ), .Y(
        XOR2_55_Y));
    AND2 AND2_24 (.A(XOR2_76_Y), .B(XOR2_7_Y), .Y(AND2_24_Y));
    AO1 AO1_40 (.A(AND2_17_Y), .B(AO1_27_Y), .C(AO1_50_Y), .Y(AO1_40_Y)
        );
    XOR2 XOR2_72 (.A(\WBINSYNCSHIFT[9] ), .B(INV_3_Y), .Y(XOR2_72_Y));
    XNOR2 XNOR2_0 (.A(\RBINSYNCSHIFT[4] ), .B(\WBINNXTSHIFT[4] ), .Y(
        XNOR2_0_Y));
    AND2 AND2_31 (.A(AND2_58_Y), .B(AND2_11_Y), .Y(AND2_31_Y));
    DFN1C0 \DFN1C0_MEM_WADDR[10]  (.D(\WBINNXTSHIFT[10] ), .CLK(WCLOCK)
        , .CLR(WRITE_RESET_P), .Q(\MEM_WADDR[10] ));
    DFN1C0 DFN1C0_15 (.D(VCC), .CLK(WCLOCK), .CLR(RESET_POLA), .Q(
        DFN1C0_15_Q));
    AO1 AO1_34 (.A(AND2_65_Y), .B(AO1_7_Y), .C(AO1_8_Y), .Y(AO1_34_Y));
    XNOR3 XNOR3_42 (.A(\RGRYSYNC[9] ), .B(\RGRYSYNC[8] ), .C(
        \RGRYSYNC[7] ), .Y(XNOR3_42_Y));
    DFN1C0 DFN1C0_12 (.D(\WGRY[11] ), .CLK(RCLOCK), .CLR(READ_RESET_P), 
        .Q(DFN1C0_12_Q));
    XOR2 \XOR2_RBINNXTSHIFT[12]  (.A(XOR2_98_Y), .B(AO1_49_Y), .Y(
        \RBINNXTSHIFT[12] ));
    XOR2 XOR2_18 (.A(\RBINNXTSHIFT[0] ), .B(\RBINNXTSHIFT[1] ), .Y(
        XOR2_18_Y));
    XNOR3 XNOR3_19 (.A(\RGRYSYNC[6] ), .B(\RGRYSYNC[5] ), .C(
        \RGRYSYNC[4] ), .Y(XNOR3_19_Y));
    DFN1C0 \DFN1C0_RGRY[11]  (.D(XOR2_6_Y), .CLK(RCLOCK), .CLR(
        READ_RESET_P), .Q(\RGRY[11] ));
    DFN1C0 \DFN1C0_WGRYSYNC[9]  (.D(DFN1C0_22_Q), .CLK(RCLOCK), .CLR(
        READ_RESET_P), .Q(\WGRYSYNC[9] ));
    XOR2 \XOR2_RBINNXTSHIFT[4]  (.A(XOR2_96_Y), .B(AO1_12_Y), .Y(
        \RBINNXTSHIFT[4] ));
    XOR2 XOR2_89 (.A(\WBINSYNCSHIFT[1] ), .B(INV_0_Y), .Y(XOR2_89_Y));
    AO1 AO1_46 (.A(XOR2_95_Y), .B(AO1_49_Y), .C(AND2_84_Y), .Y(
        AO1_46_Y));
    DFN1C0 \DFN1C0_MEM_WADDR[8]  (.D(\WBINNXTSHIFT[8] ), .CLK(WCLOCK), 
        .CLR(WRITE_RESET_P), .Q(\MEM_WADDR[8] ));
    XNOR3 XNOR3_22 (.A(\WGRYSYNC[12] ), .B(\WGRYSYNC[11] ), .C(
        \WGRYSYNC[10] ), .Y(XNOR3_22_Y));
    DFN1C0 \DFN1C0_RGRY[1]  (.D(XOR2_28_Y), .CLK(RCLOCK), .CLR(
        READ_RESET_P), .Q(\RGRY[1] ));
    DFN1C0 \DFN1C0_RGRYSYNC[5]  (.D(DFN1C0_14_Q), .CLK(WCLOCK), .CLR(
        WRITE_RESET_P), .Q(\RGRYSYNC[5] ));
    DFN1C0 \DFN1C0_WGRY[3]  (.D(XOR2_73_Y), .CLK(WCLOCK), .CLR(
        WRITE_RESET_P), .Q(\WGRY[3] ));
    XOR2 XOR2_8 (.A(\MEM_RADDR[11] ), .B(GND), .Y(XOR2_8_Y));
    XOR2 \XOR2_RBINNXTSHIFT[6]  (.A(XOR2_88_Y), .B(AO1_6_Y), .Y(
        \RBINNXTSHIFT[6] ));
    AO1 AO1_43 (.A(AND2_42_Y), .B(AO1_44_Y), .C(AO1_11_Y), .Y(AO1_43_Y)
        );
    XNOR3 XNOR3_39 (.A(\RGRYSYNC[6] ), .B(\RGRYSYNC[5] ), .C(
        \RGRYSYNC[4] ), .Y(XNOR3_39_Y));
    XOR2 XOR2_30 (.A(\MEM_WADDR[11] ), .B(GND), .Y(XOR2_30_Y));
    XOR2 \XOR2_RDIFF[0]  (.A(\WBINSYNCSHIFT[0] ), .B(\RBINNXTSHIFT[0] )
        , .Y(\RDIFF[0] ));
    AND2 AND2_38 (.A(\MEM_RADDR[10] ), .B(GND), .Y(AND2_38_Y));
    AND2 AND2_35 (.A(\WBINSYNCSHIFT[11] ), .B(INV_8_Y), .Y(AND2_35_Y));
    INV MEMREBUBBLE (.A(MEMORYRE), .Y(MEMRENEG));
    XNOR2 \XNOR2_RDIFF[1]  (.A(XOR2_89_Y), .B(NOR2A_0_Y), .Y(
        \RDIFF[1] ));
    DFN1C0 \DFN1C0_MEM_WADDR[7]  (.D(\WBINNXTSHIFT[7] ), .CLK(WCLOCK), 
        .CLR(WRITE_RESET_P), .Q(\MEM_WADDR[7] ));
    DFN1C0 \DFN1C0_WGRY[11]  (.D(XOR2_3_Y), .CLK(WCLOCK), .CLR(
        WRITE_RESET_P), .Q(\WGRY[11] ));
    AND2 AND2_29 (.A(AND2_58_Y), .B(AND2_64_Y), .Y(AND2_29_Y));
    DFN1C0 \DFN1C0_MEM_RADDR[4]  (.D(\RBINNXTSHIFT[4] ), .CLK(RCLOCK), 
        .CLR(READ_RESET_P), .Q(\MEM_RADDR[4] ));
    XNOR3 XNOR3_7 (.A(\RGRYSYNC[9] ), .B(\RGRYSYNC[8] ), .C(
        \RGRYSYNC[7] ), .Y(XNOR3_7_Y));
    XNOR3 XNOR3_46 (.A(\RGRYSYNC[12] ), .B(\RGRYSYNC[11] ), .C(
        \RGRYSYNC[10] ), .Y(XNOR3_46_Y));
    XOR2 \XOR2_WBINNXTSHIFT[12]  (.A(XOR2_17_Y), .B(AO1_22_Y), .Y(
        \WBINNXTSHIFT[12] ));
    XOR2 XOR2_34 (.A(\MEM_WADDR[12] ), .B(GND), .Y(XOR2_34_Y));
    XOR2 XOR2_31 (.A(\MEM_RADDR[5] ), .B(GND), .Y(XOR2_31_Y));
    AND2 AND2_3 (.A(\MEM_WADDR[10] ), .B(GND), .Y(AND2_3_Y));
    DFN1C0 \DFN1C0_MEM_WADDR[11]  (.D(\WBINNXTSHIFT[11] ), .CLK(WCLOCK)
        , .CLR(WRITE_RESET_P), .Q(\MEM_WADDR[11] ));
    AO1 AO1_49 (.A(AND2_83_Y), .B(AO1_29_Y), .C(AO1_0_Y), .Y(AO1_49_Y));
    AND2 AND2_30 (.A(XOR2_41_Y), .B(XOR2_94_Y), .Y(AND2_30_Y));
    XOR2 \XOR2_WBINNXTSHIFT[4]  (.A(XOR2_99_Y), .B(AO1_36_Y), .Y(
        \WBINNXTSHIFT[4] ));
    XNOR3 XNOR3_26 (.A(\WGRYSYNC[9] ), .B(\WGRYSYNC[8] ), .C(
        \WGRYSYNC[7] ), .Y(XNOR3_26_Y));
    XNOR2 XNOR2_6 (.A(\RBINSYNCSHIFT[10] ), .B(\WBINNXTSHIFT[10] ), .Y(
        XNOR2_6_Y));
    INV RESETBUBBLE (.A(RESET), .Y(RESET_POLA));
    AND2 AND2_14 (.A(\MEM_WADDR[5] ), .B(GND), .Y(AND2_14_Y));
    INV INV_4 (.A(NOR2A_0_Y), .Y(INV_4_Y));
    AND2 AND2_74 (.A(\WBINSYNCSHIFT[7] ), .B(INV_7_Y), .Y(AND2_74_Y));
    XOR2 XOR2_77 (.A(\MEM_WADDR[5] ), .B(GND), .Y(XOR2_77_Y));
    AND2 AND2_32 (.A(AND2_15_Y), .B(XOR2_41_Y), .Y(AND2_32_Y));
    XOR2 \XOR2_WBINNXTSHIFT[6]  (.A(XOR2_78_Y), .B(AO1_17_Y), .Y(
        \WBINNXTSHIFT[6] ));
    DFN1C0 \DFN1C0_MEM_RADDR[5]  (.D(\RBINNXTSHIFT[5] ), .CLK(RCLOCK), 
        .CLR(READ_RESET_P), .Q(\MEM_RADDR[5] ));
    AND3 AND3_8 (.A(AND3_9_Y), .B(AND3_7_Y), .C(AND3_6_Y), .Y(AND3_8_Y)
        );
    XOR3 XOR3_4 (.A(\WGRYSYNC[12] ), .B(\WGRYSYNC[11] ), .C(
        \WGRYSYNC[10] ), .Y(XOR3_4_Y));
    XOR2 XOR2_46 (.A(\MEM_RADDR[2] ), .B(GND), .Y(XOR2_46_Y));
    XNOR2 XNOR2_11 (.A(\RBINSYNCSHIFT[11] ), .B(\WBINNXTSHIFT[11] ), 
        .Y(XNOR2_11_Y));
    AO1 AO1_2 (.A(AND2_21_Y), .B(AO1_4_Y), .C(AO1_10_Y), .Y(AO1_2_Y));
    DFN1C0 \DFN1C0_MEM_RADDR[8]  (.D(\RBINNXTSHIFT[8] ), .CLK(RCLOCK), 
        .CLR(READ_RESET_P), .Q(\MEM_RADDR[8] ));
    DFN1C0 \DFN1C0_WGRY[0]  (.D(XOR2_42_Y), .CLK(WCLOCK), .CLR(
        WRITE_RESET_P), .Q(\WGRY[0] ));
    DFN1C0 \DFN1C0_RDCNT[7]  (.D(\RDIFF[7] ), .CLK(RCLOCK), .CLR(
        READ_RESET_P), .Q(RDCNT[7]));
    XOR2 XOR2_75 (.A(\RBINNXTSHIFT[6] ), .B(\RBINNXTSHIFT[7] ), .Y(
        XOR2_75_Y));
    AND2 AND2_26 (.A(AND2_31_Y), .B(XOR2_79_Y), .Y(AND2_26_Y));
    XOR2 XOR2_99 (.A(\MEM_WADDR[4] ), .B(GND), .Y(XOR2_99_Y));
    XOR2 XOR2_9 (.A(\MEM_RADDR[9] ), .B(GND), .Y(XOR2_9_Y));
    AND3 AND3_5 (.A(XNOR2_1_Y), .B(XNOR2_17_Y), .C(XNOR2_21_Y), .Y(
        AND3_5_Y));
    XNOR2 \XNOR2_WBINSYNCSHIFT[5]  (.A(XNOR3_14_Y), .B(XNOR3_33_Y), .Y(
        \WBINSYNCSHIFT[5] ));
    INV INV_12 (.A(\RBINNXTSHIFT[4] ), .Y(INV_12_Y));
    XOR2 XOR2_59 (.A(\WBINNXTSHIFT[7] ), .B(\WBINNXTSHIFT[8] ), .Y(
        XOR2_59_Y));
    AND2 AND2_23 (.A(AND2_12_Y), .B(XOR2_0_Y), .Y(AND2_23_Y));
    DFN1C0 \DFN1C0_MEM_WADDR[9]  (.D(\WBINNXTSHIFT[9] ), .CLK(WCLOCK), 
        .CLR(WRITE_RESET_P), .Q(\MEM_WADDR[9] ));
    DFN1C0 \DFN1C0_WGRYSYNC[1]  (.D(DFN1C0_10_Q), .CLK(RCLOCK), .CLR(
        READ_RESET_P), .Q(\WGRYSYNC[1] ));
    XNOR2 XNOR2_4 (.A(\RBINNXTSHIFT[11] ), .B(\WBINSYNCSHIFT[11] ), .Y(
        XNOR2_4_Y));
    DFN1C0 \DFN1C0_RGRY[8]  (.D(XOR2_74_Y), .CLK(RCLOCK), .CLR(
        READ_RESET_P), .Q(\RGRY[8] ));
    XOR2 XOR2_5 (.A(\MEM_RADDR[7] ), .B(GND), .Y(XOR2_5_Y));
    XNOR3 XNOR3_47 (.A(\RGRYSYNC[3] ), .B(XOR3_2_Y), .C(XNOR3_1_Y), .Y(
        XNOR3_47_Y));
    XNOR2 XNOR2_20 (.A(\RBINNXTSHIFT[7] ), .B(\WBINSYNCSHIFT[7] ), .Y(
        XNOR2_20_Y));
    DFN1C0 DFN1C0_16 (.D(\RGRY[7] ), .CLK(WCLOCK), .CLR(WRITE_RESET_P), 
        .Q(DFN1C0_16_Q));
    XNOR3 XNOR3_11 (.A(\WGRYSYNC[0] ), .B(XNOR3_35_Y), .C(XNOR3_48_Y), 
        .Y(XNOR3_11_Y));
    AO1 AO1_28 (.A(AND2_8_Y), .B(AO1_2_Y), .C(AO1_23_Y), .Y(AO1_28_Y));
    AND2 AND2_19 (.A(\MEM_RADDR[5] ), .B(GND), .Y(AND2_19_Y));
    DFN1C0 DFN1C0_6 (.D(\RGRY[2] ), .CLK(WCLOCK), .CLR(WRITE_RESET_P), 
        .Q(DFN1C0_6_Q));
    AND2 AND2_79 (.A(XOR2_13_Y), .B(XOR2_4_Y), .Y(AND2_79_Y));
    XNOR2 \XNOR2_WBINSYNCSHIFT[7]  (.A(XOR3_6_Y), .B(XNOR3_25_Y), .Y(
        \WBINSYNCSHIFT[7] ));
    DFN1C0 \DFN1C0_MEM_RADDR[6]  (.D(\RBINNXTSHIFT[6] ), .CLK(RCLOCK), 
        .CLR(READ_RESET_P), .Q(\MEM_RADDR[6] ));
    XOR2 XOR2_86 (.A(\MEM_WADDR[3] ), .B(GND), .Y(XOR2_86_Y));
    XNOR3 XNOR3_27 (.A(\WGRYSYNC[9] ), .B(\WGRYSYNC[8] ), .C(
        \WGRYSYNC[7] ), .Y(XNOR3_27_Y));
    XOR2 XOR2_22 (.A(\MEM_WADDR[2] ), .B(GND), .Y(XOR2_22_Y));
    DFN1C0 \DFN1C0_RDCNT[1]  (.D(\RDIFF[1] ), .CLK(RCLOCK), .CLR(
        READ_RESET_P), .Q(RDCNT[1]));
    RAM4K9 RAM4K9_QXI (.ADDRA11(\MEM_WADDR[11] ), .ADDRA10(
        \MEM_WADDR[10] ), .ADDRA9(\MEM_WADDR[9] ), .ADDRA8(
        \MEM_WADDR[8] ), .ADDRA7(\MEM_WADDR[7] ), .ADDRA6(
        \MEM_WADDR[6] ), .ADDRA5(\MEM_WADDR[5] ), .ADDRA4(
        \MEM_WADDR[4] ), .ADDRA3(\MEM_WADDR[3] ), .ADDRA2(
        \MEM_WADDR[2] ), .ADDRA1(\MEM_WADDR[1] ), .ADDRA0(
        \MEM_WADDR[0] ), .ADDRB11(\MEM_RADDR[11] ), .ADDRB10(
        \MEM_RADDR[10] ), .ADDRB9(\MEM_RADDR[9] ), .ADDRB8(
        \MEM_RADDR[8] ), .ADDRB7(\MEM_RADDR[7] ), .ADDRB6(
        \MEM_RADDR[6] ), .ADDRB5(\MEM_RADDR[5] ), .ADDRB4(
        \MEM_RADDR[4] ), .ADDRB3(\MEM_RADDR[3] ), .ADDRB2(
        \MEM_RADDR[2] ), .ADDRB1(\MEM_RADDR[1] ), .ADDRB0(
        \MEM_RADDR[0] ), .DINA8(GND), .DINA7(GND), .DINA6(GND), .DINA5(
        GND), .DINA4(GND), .DINA3(GND), .DINA2(GND), .DINA1(GND), 
        .DINA0(DATA), .DINB8(GND), .DINB7(GND), .DINB6(GND), .DINB5(
        GND), .DINB4(GND), .DINB3(GND), .DINB2(GND), .DINB1(GND), 
        .DINB0(GND), .WIDTHA0(GND), .WIDTHA1(GND), .WIDTHB0(GND), 
        .WIDTHB1(GND), .PIPEA(GND), .PIPEB(GND), .WMODEA(GND), .WMODEB(
        GND), .BLKA(MEMWENEG), .BLKB(MEMRENEG), .WENA(GND), .WENB(VCC), 
        .CLKA(WCLOCK), .CLKB(RCLOCK), .RESET(WRITE_RESET_P), .DOUTA8(), 
        .DOUTA7(), .DOUTA6(), .DOUTA5(), .DOUTA4(), .DOUTA3(), .DOUTA2(
        ), .DOUTA1(), .DOUTA0(RAM4K9_QXI_DOUTA0), .DOUTB8(), .DOUTB7(), 
        .DOUTB6(), .DOUTB5(), .DOUTB4(), .DOUTB3(), .DOUTB2(), .DOUTB1(
        ), .DOUTB0(QXI));
    XNOR3 \XNOR3_RBINSYNCSHIFT[8]  (.A(\RGRYSYNC[9] ), .B(
        \RGRYSYNC[8] ), .C(XNOR3_24_Y), .Y(\RBINSYNCSHIFT[8] ));
    AO1 AO1_1 (.A(XOR2_40_Y), .B(AND2_39_Y), .C(AND2_66_Y), .Y(AO1_1_Y)
        );
    XOR2 \XOR2_RDIFF[9]  (.A(XOR2_72_Y), .B(AO1_5_Y), .Y(\RDIFF[9] ));
    DFN1C0 DFN1C0_10 (.D(\WGRY[1] ), .CLK(RCLOCK), .CLR(READ_RESET_P), 
        .Q(DFN1C0_10_Q));
    XOR2 XOR2_13 (.A(\MEM_RADDR[2] ), .B(GND), .Y(XOR2_13_Y));
    DFN1C0 \DFN1C0_WGRYSYNC[2]  (.D(DFN1C0_11_Q), .CLK(RCLOCK), .CLR(
        READ_RESET_P), .Q(\WGRYSYNC[2] ));
    XNOR3 XNOR3_31 (.A(\WGRYSYNC[9] ), .B(\WGRYSYNC[8] ), .C(
        \WGRYSYNC[7] ), .Y(XNOR3_31_Y));
    INV INV_6 (.A(\RBINNXTSHIFT[12] ), .Y(INV_6_Y));
    DFN1C0 \DFN1C0_WGRYSYNC[0]  (.D(DFN1C0_13_Q), .CLK(RCLOCK), .CLR(
        READ_RESET_P), .Q(\WGRYSYNC[0] ));
    XNOR2 XNOR2_18 (.A(\RBINNXTSHIFT[6] ), .B(\WBINSYNCSHIFT[6] ), .Y(
        XNOR2_18_Y));
    AND2 AND2_51 (.A(\WBINSYNCSHIFT[4] ), .B(INV_12_Y), .Y(AND2_51_Y));
    AO1 AO1_3 (.A(XOR2_26_Y), .B(AO1_41_Y), .C(AND2_35_Y), .Y(AO1_3_Y));
    AND2 AND2_64 (.A(AND2_11_Y), .B(AND2_17_Y), .Y(AND2_64_Y));
    AND2 AND2_47 (.A(AND2_87_Y), .B(XOR2_15_Y), .Y(AND2_47_Y));
    AO1 AO1_51 (.A(XOR2_14_Y), .B(AO1_5_Y), .C(AND2_60_Y), .Y(AO1_51_Y)
        );
    XNOR3 XNOR3_44 (.A(\RGRYSYNC[6] ), .B(\RGRYSYNC[5] ), .C(
        \RGRYSYNC[4] ), .Y(XNOR3_44_Y));
    AO1 AO1_18 (.A(XOR2_1_Y), .B(AO1_17_Y), .C(AND2_78_Y), .Y(AO1_18_Y)
        );
    XOR2 XOR2_48 (.A(\WBINSYNCSHIFT[10] ), .B(INV_11_Y), .Y(XOR2_48_Y));
    AO1 AO1_47 (.A(XOR2_85_Y), .B(AND2_34_Y), .C(AND2_46_Y), .Y(
        AO1_47_Y));
    XOR2 \XOR2_RBINNXTSHIFT[3]  (.A(XOR2_69_Y), .B(AO1_35_Y), .Y(
        \RBINNXTSHIFT[3] ));
    DFN1C0 DFN1C0_3 (.D(VCC), .CLK(RCLOCK), .CLR(RESET_POLA), .Q(
        DFN1C0_3_Q));
    DFN1C0 \DFN1C0_MEM_RADDR[7]  (.D(\RBINNXTSHIFT[7] ), .CLK(RCLOCK), 
        .CLR(READ_RESET_P), .Q(\MEM_RADDR[7] ));
    AND2 AND2_16 (.A(AND2_24_Y), .B(XOR2_13_Y), .Y(AND2_16_Y));
    XNOR3 XNOR3_18 (.A(\WGRYSYNC[3] ), .B(XOR3_0_Y), .C(XNOR3_27_Y), 
        .Y(XNOR3_18_Y));
    XOR2 \XOR2_RDIFF[8]  (.A(XOR2_60_Y), .B(AO1_14_Y), .Y(\RDIFF[8] ));
    XNOR3 XNOR3_24 (.A(\RGRYSYNC[12] ), .B(\RGRYSYNC[11] ), .C(
        \RGRYSYNC[10] ), .Y(XNOR3_24_Y));
    AND2 AND2_76 (.A(AND2_58_Y), .B(XOR2_25_Y), .Y(AND2_76_Y));
    AO1 AO1_38 (.A(AND2_63_Y), .B(AO1_5_Y), .C(AO1_43_Y), .Y(AO1_38_Y));
    DFN1C0 \DFN1C0_WGRY[9]  (.D(XOR2_21_Y), .CLK(WCLOCK), .CLR(
        WRITE_RESET_P), .Q(\WGRY[9] ));
    XOR2 XOR2_62 (.A(\WBINNXTSHIFT[8] ), .B(\WBINNXTSHIFT[9] ), .Y(
        XOR2_62_Y));
    AND2 AND2_13 (.A(\MEM_WADDR[2] ), .B(GND), .Y(AND2_13_Y));
    AND2 AND2_87 (.A(AND2_24_Y), .B(AND2_79_Y), .Y(AND2_87_Y));
    DFN1C0 DFN1C0_18 (.D(\RGRY[3] ), .CLK(WCLOCK), .CLR(WRITE_RESET_P), 
        .Q(DFN1C0_18_Q));
    AND2 AND2_73 (.A(\MEM_WADDR[9] ), .B(GND), .Y(AND2_73_Y));
    XOR2 XOR2_10 (.A(\WBINSYNCSHIFT[1] ), .B(INV_0_Y), .Y(XOR2_10_Y));
    XNOR2 XNOR2_1 (.A(\RBINSYNCSHIFT[0] ), .B(\WBINNXTSHIFT[0] ), .Y(
        XNOR2_1_Y));
    XNOR3 XNOR3_38 (.A(\WGRYSYNC[6] ), .B(\WGRYSYNC[5] ), .C(
        \WGRYSYNC[4] ), .Y(XNOR3_38_Y));
    AND2 AND2_58 (.A(AND2_41_Y), .B(AND2_36_Y), .Y(AND2_58_Y));
    AND2 AND2_55 (.A(\WBINSYNCSHIFT[2] ), .B(INV_9_Y), .Y(AND2_55_Y));
    INV INV_8 (.A(\RBINNXTSHIFT[11] ), .Y(INV_8_Y));
    XNOR3 XNOR3_6 (.A(\RGRYSYNC[12] ), .B(\RGRYSYNC[11] ), .C(
        \RGRYSYNC[10] ), .Y(XNOR3_6_Y));
    DFN1C0 \DFN1C0_RDCNT[8]  (.D(\RDIFF[8] ), .CLK(RCLOCK), .CLR(
        READ_RESET_P), .Q(RDCNT[8]));
    DFN1C0 \DFN1C0_RGRY[4]  (.D(XOR2_84_Y), .CLK(RCLOCK), .CLR(
        READ_RESET_P), .Q(\RGRY[4] ));
    DFN1C0 DFN1C0_2 (.D(\WGRY[10] ), .CLK(RCLOCK), .CLR(READ_RESET_P), 
        .Q(DFN1C0_2_Q));
    XOR2 XOR2_88 (.A(\MEM_RADDR[6] ), .B(GND), .Y(XOR2_88_Y));
    XNOR3 XNOR3_43 (.A(\RGRYSYNC[6] ), .B(\RGRYSYNC[5] ), .C(
        \RGRYSYNC[4] ), .Y(XNOR3_43_Y));
    XOR2 XOR2_96 (.A(\MEM_RADDR[4] ), .B(GND), .Y(XOR2_96_Y));
    AND2 AND2_69 (.A(AND2_94_Y), .B(XOR2_95_Y), .Y(AND2_69_Y));
    DFN1C0 \DFN1C0_MEM_WADDR[2]  (.D(\WBINNXTSHIFT[2] ), .CLK(WCLOCK), 
        .CLR(WRITE_RESET_P), .Q(\MEM_WADDR[2] ));
    XOR2 XOR2_79 (.A(\MEM_WADDR[10] ), .B(GND), .Y(XOR2_79_Y));
    XOR3 XOR3_3 (.A(\WGRYSYNC[12] ), .B(\WGRYSYNC[11] ), .C(
        \WGRYSYNC[10] ), .Y(XOR3_3_Y));
    XOR2 XOR2_27 (.A(\MEM_RADDR[5] ), .B(GND), .Y(XOR2_27_Y));
    AND2 AND2_MEMORYRE (.A(NAND2_1_Y), .B(RE), .Y(MEMORYRE));
    XOR2 \XOR2_WBINNXTSHIFT[3]  (.A(XOR2_90_Y), .B(AO1_37_Y), .Y(
        \WBINNXTSHIFT[3] ));
    XOR2 XOR2_7 (.A(\MEM_RADDR[1] ), .B(GND), .Y(XOR2_7_Y));
    AND2 AND2_5 (.A(\MEM_RADDR[4] ), .B(GND), .Y(AND2_5_Y));
    XOR2 XOR2_56 (.A(\MEM_WADDR[9] ), .B(GND), .Y(XOR2_56_Y));
    XOR2 XOR2_14 (.A(\WBINSYNCSHIFT[9] ), .B(INV_3_Y), .Y(XOR2_14_Y));
    AND2 AND2_91 (.A(\MEM_RADDR[0] ), .B(MEMORYRE), .Y(AND2_91_Y));
    AND2 AND2_50 (.A(\WBINSYNCSHIFT[8] ), .B(INV_1_Y), .Y(AND2_50_Y));
    XNOR3 XNOR3_23 (.A(\RGRYSYNC[9] ), .B(\RGRYSYNC[8] ), .C(
        \RGRYSYNC[7] ), .Y(XNOR3_23_Y));
    XNOR3 XNOR3_1 (.A(\RGRYSYNC[9] ), .B(\RGRYSYNC[8] ), .C(
        \RGRYSYNC[7] ), .Y(XNOR3_1_Y));
    DFN1C0 DFN1C0_7 (.D(\RGRY[10] ), .CLK(WCLOCK), .CLR(WRITE_RESET_P), 
        .Q(DFN1C0_7_Q));
    XNOR2 XNOR2_3 (.A(\RBINSYNCSHIFT[9] ), .B(\WBINNXTSHIFT[9] ), .Y(
        XNOR2_3_Y));
    XOR2 XOR2_11 (.A(\WBINSYNCSHIFT[2] ), .B(INV_9_Y), .Y(XOR2_11_Y));
    XNOR2 XNOR2_22 (.A(\RBINNXTSHIFT[12] ), .B(READDOMAIN_WMSB), .Y(
        XNOR2_22_Y));
    XOR3 XOR3_6 (.A(\WGRYSYNC[12] ), .B(\WGRYSYNC[11] ), .C(
        \WGRYSYNC[10] ), .Y(XOR3_6_Y));
    AND2 AND2_52 (.A(AND2_87_Y), .B(AND2_27_Y), .Y(AND2_52_Y));
    XOR2 XOR2_25 (.A(\MEM_WADDR[8] ), .B(GND), .Y(XOR2_25_Y));
    XNOR2 XNOR2_15 (.A(\RBINSYNCSHIFT[6] ), .B(\WBINNXTSHIFT[6] ), .Y(
        XNOR2_15_Y));
    AO1 AO1_22 (.A(AND2_64_Y), .B(AO1_9_Y), .C(AO1_40_Y), .Y(AO1_22_Y));
    XNOR3 XNOR3_3 (.A(\RGRYSYNC[9] ), .B(\RGRYSYNC[8] ), .C(
        \RGRYSYNC[7] ), .Y(XNOR3_3_Y));
    XNOR2 \XNOR2_RBINSYNCSHIFT[7]  (.A(XOR3_1_Y), .B(XNOR3_51_Y), .Y(
        \RBINSYNCSHIFT[7] ));
    DFN1C0 \DFN1C0_RGRYSYNC[10]  (.D(DFN1C0_7_Q), .CLK(WCLOCK), .CLR(
        WRITE_RESET_P), .Q(\RGRYSYNC[10] ));
    AO1 AO1_55 (.A(XOR2_5_Y), .B(AND2_1_Y), .C(AND2_43_Y), .Y(AO1_55_Y)
        );
    DFN1C0 \DFN1C0_RGRYSYNC[9]  (.D(DFN1C0_1_Q), .CLK(WCLOCK), .CLR(
        WRITE_RESET_P), .Q(\RGRYSYNC[9] ));
    AND2 AND2_34 (.A(\MEM_RADDR[8] ), .B(GND), .Y(AND2_34_Y));
    AO1 AO1_41 (.A(AND2_88_Y), .B(AO1_5_Y), .C(AO1_44_Y), .Y(AO1_41_Y));
    AND2 AND2_66 (.A(\MEM_WADDR[1] ), .B(GND), .Y(AND2_66_Y));
    AO1 AO1_6 (.A(AND2_27_Y), .B(AO1_12_Y), .C(AO1_16_Y), .Y(AO1_6_Y));
    XNOR3 XNOR3_15 (.A(\WGRYSYNC[6] ), .B(\WGRYSYNC[5] ), .C(
        \WGRYSYNC[4] ), .Y(XNOR3_15_Y));
    AND2 AND2_95 (.A(AND2_0_Y), .B(AND2_70_Y), .Y(AND2_95_Y));
    DFN1C0 \DFN1C0_MEM_RADDR[3]  (.D(\RBINNXTSHIFT[3] ), .CLK(RCLOCK), 
        .CLR(READ_RESET_P), .Q(\MEM_RADDR[3] ));
    XOR2 XOR2_67 (.A(\MEM_WADDR[11] ), .B(GND), .Y(XOR2_67_Y));
    DFN1C0 DFN1C0_23 (.D(\WGRY[8] ), .CLK(RCLOCK), .CLR(READ_RESET_P), 
        .Q(DFN1C0_23_Q));
    AND2 AND2_63 (.A(AND2_88_Y), .B(AND2_42_Y), .Y(AND2_63_Y));
    AND3 AND3_2 (.A(AND3_4_Y), .B(AND3_5_Y), .C(AND3_3_Y), .Y(AND3_2_Y)
        );
    DFN1E1C0 DFN1E1C0_Q (.D(QXI), .CLK(RCLOCK), .CLR(READ_RESET_P), .E(
        DVLDI), .Q(Q));
    AO1 AO1_12 (.A(AND2_79_Y), .B(AO1_24_Y), .C(AO1_45_Y), .Y(AO1_12_Y)
        );
    XOR2 XOR2_32 (.A(\WBINSYNCSHIFT[2] ), .B(INV_9_Y), .Y(XOR2_32_Y));
    OR3 OR3_0 (.A(AND2_37_Y), .B(AND2_22_Y), .C(AND2_67_Y), .Y(OR3_0_Y)
        );
    XOR2 XOR2_98 (.A(\MEM_RADDR[12] ), .B(GND), .Y(XOR2_98_Y));
    XNOR3 XNOR3_35 (.A(\WGRYSYNC[12] ), .B(\WGRYSYNC[11] ), .C(
        \WGRYSYNC[10] ), .Y(XNOR3_35_Y));
    XOR2 \XOR2_RDIFF[7]  (.A(XOR2_38_Y), .B(AO1_28_Y), .Y(\RDIFF[7] ));
    AND2 AND2_9 (.A(\MEM_WADDR[3] ), .B(GND), .Y(AND2_9_Y));
    XOR2 XOR2_65 (.A(\MEM_WADDR[7] ), .B(GND), .Y(XOR2_65_Y));
    AND2 AND2_90 (.A(\WBINSYNCSHIFT[6] ), .B(INV_5_Y), .Y(AND2_90_Y));
    XOR2 XOR2_58 (.A(\RBINNXTSHIFT[3] ), .B(\RBINNXTSHIFT[4] ), .Y(
        XOR2_58_Y));
    XOR2 XOR2_43 (.A(\RBINNXTSHIFT[9] ), .B(\RBINNXTSHIFT[10] ), .Y(
        XOR2_43_Y));
    XOR2 \XOR2_RDIFF[2]  (.A(XOR2_32_Y), .B(OR3_0_Y), .Y(\RDIFF[2] ));
    AO1 AO1_32 (.A(XOR2_71_Y), .B(AO1_6_Y), .C(AND2_1_Y), .Y(AO1_32_Y));
    INV INV_2 (.A(\RBINNXTSHIFT[3] ), .Y(INV_2_Y));
    XNOR2 \XNOR2_RBINSYNCSHIFT[3]  (.A(XNOR3_39_Y), .B(XNOR3_47_Y), .Y(
        \RBINSYNCSHIFT[3] ));
    AND2 AND2_92 (.A(\WBINSYNCSHIFT[3] ), .B(INV_2_Y), .Y(AND2_92_Y));
    DFN1C0 \DFN1C0_RGRYSYNC[12]  (.D(DFN1C0_19_Q), .CLK(WCLOCK), .CLR(
        WRITE_RESET_P), .Q(\RGRYSYNC[12] ));
    AO1 AO1_9 (.A(AND2_36_Y), .B(AO1_36_Y), .C(AO1_34_Y), .Y(AO1_9_Y));
    XOR2 \XOR2_RDIFF[12]  (.A(XOR2_61_Y), .B(AO1_3_Y), .Y(\RDIFF[12] ));
    DFN1C0 DFN1C0_DVLDX (.D(DVLDI), .CLK(RCLOCK), .CLR(READ_RESET_P), 
        .Q(DVLDX));
    NAND2 NAND2_0 (.A(FULL), .B(VCC), .Y(NAND2_0_Y));
    AND2 AND2_39 (.A(\MEM_WADDR[0] ), .B(MEMORYWE), .Y(AND2_39_Y));
    XNOR3 XNOR3_0 (.A(\RGRYSYNC[9] ), .B(\RGRYSYNC[8] ), .C(
        \RGRYSYNC[7] ), .Y(XNOR3_0_Y));
    DFN1C0 \DFN1C0_WGRYSYNC[10]  (.D(DFN1C0_2_Q), .CLK(RCLOCK), .CLR(
        READ_RESET_P), .Q(\WGRYSYNC[10] ));
    DFN1C0 \DFN1C0_RGRY[6]  (.D(XOR2_75_Y), .CLK(RCLOCK), .CLR(
        READ_RESET_P), .Q(\RGRY[6] ));
    XOR2 XOR2_76 (.A(\MEM_RADDR[0] ), .B(MEMORYRE), .Y(XOR2_76_Y));
    AND2 AND2_27 (.A(XOR2_15_Y), .B(XOR2_31_Y), .Y(AND2_27_Y));
    DFN1C0 DFN1C0_DVLDI (.D(AND2A_0_Y), .CLK(RCLOCK), .CLR(
        READ_RESET_P), .Q(DVLDI));
    XNOR2 XNOR2_10 (.A(\RBINNXTSHIFT[5] ), .B(\WBINSYNCSHIFT[5] ), .Y(
        XNOR2_10_Y));
    AO1 AO1_54 (.A(XOR2_68_Y), .B(AO1_26_Y), .C(AND2_38_Y), .Y(
        AO1_54_Y));
    AND2 AND2_MEMORYWE (.A(NAND2_0_Y), .B(WE), .Y(MEMORYWE));
    XOR2 XOR2_83 (.A(\MEM_RADDR[7] ), .B(GND), .Y(XOR2_83_Y));
    AO1 AO1_20 (.A(XOR2_15_Y), .B(AO1_12_Y), .C(AND2_5_Y), .Y(AO1_20_Y)
        );
    DFN1C0 \DFN1C0_WGRY[2]  (.D(XOR2_23_Y), .CLK(WCLOCK), .CLR(
        WRITE_RESET_P), .Q(\WGRY[2] ));
    AO1 AO1_0 (.A(AND2_61_Y), .B(AO1_47_Y), .C(AO1_25_Y), .Y(AO1_0_Y));
    XOR2 XOR2_29 (.A(\WBINSYNCSHIFT[5] ), .B(INV_10_Y), .Y(XOR2_29_Y));
    DFN1C0 \DFN1C0_WGRYSYNC[8]  (.D(DFN1C0_23_Q), .CLK(RCLOCK), .CLR(
        READ_RESET_P), .Q(\WGRYSYNC[8] ));
    AO1 AO1_45 (.A(XOR2_4_Y), .B(AND2_20_Y), .C(AND2_68_Y), .Y(
        AO1_45_Y));
    XOR2 XOR2_40 (.A(\MEM_WADDR[1] ), .B(GND), .Y(XOR2_40_Y));
    DFN1C0 \DFN1C0_RGRYSYNC[1]  (.D(DFN1C0_0_Q), .CLK(WCLOCK), .CLR(
        WRITE_RESET_P), .Q(\RGRYSYNC[1] ));
    XOR3 XOR3_0 (.A(\WGRYSYNC[12] ), .B(\WGRYSYNC[11] ), .C(
        \WGRYSYNC[10] ), .Y(XOR3_0_Y));
    XOR2 XOR2_2 (.A(\MEM_WADDR[8] ), .B(GND), .Y(XOR2_2_Y));
    DFN1C0 DFN1C0_8 (.D(\WGRY[7] ), .CLK(RCLOCK), .CLR(READ_RESET_P), 
        .Q(DFN1C0_8_Q));
    DFN1C0 \DFN1C0_RGRY[5]  (.D(XOR2_92_Y), .CLK(RCLOCK), .CLR(
        READ_RESET_P), .Q(\RGRY[5] ));
    DFN1C0 \DFN1C0_RDCNT[0]  (.D(\RDIFF[0] ), .CLK(RCLOCK), .CLR(
        READ_RESET_P), .Q(RDCNT[0]));
    XNOR3 XNOR3_10 (.A(\RGRYSYNC[6] ), .B(\RGRYSYNC[5] ), .C(
        XNOR3_45_Y), .Y(XNOR3_10_Y));
    AND2A AND2A_0 (.A(EMPTY), .B(RE), .Y(AND2A_0_Y));
    XOR2 XOR2_37 (.A(\WBINNXTSHIFT[5] ), .B(\WBINNXTSHIFT[6] ), .Y(
        XOR2_37_Y));
    AND2 AND2_36 (.A(AND2_86_Y), .B(AND2_65_Y), .Y(AND2_36_Y));
    AO1 AO1_26 (.A(AND2_70_Y), .B(AO1_29_Y), .C(AO1_47_Y), .Y(AO1_26_Y)
        );
    DFN1C0 \DFN1C0_WGRY[10]  (.D(XOR2_54_Y), .CLK(WCLOCK), .CLR(
        WRITE_RESET_P), .Q(\WGRY[10] ));
    XNOR3 \XNOR3_WBINSYNCSHIFT[0]  (.A(XNOR3_15_Y), .B(XNOR3_34_Y), .C(
        XNOR3_11_Y), .Y(\WBINSYNCSHIFT[0] ));
    DFN1C0 \DFN1C0_RGRY[7]  (.D(XOR2_24_Y), .CLK(RCLOCK), .CLR(
        READ_RESET_P), .Q(\RGRY[7] ));
    AND3 AND3_9 (.A(XNOR2_18_Y), .B(XNOR2_20_Y), .C(XNOR2_16_Y), .Y(
        AND3_9_Y));
    XOR3 XOR3_5 (.A(\RGRYSYNC[12] ), .B(\RGRYSYNC[11] ), .C(
        \RGRYSYNC[10] ), .Y(XOR3_5_Y));
    XOR2 \XOR2_RBINNXTSHIFT[5]  (.A(XOR2_27_Y), .B(AO1_20_Y), .Y(
        \RBINNXTSHIFT[5] ));
    AO1 AO1_23 (.A(XOR2_44_Y), .B(AND2_53_Y), .C(AND2_90_Y), .Y(
        AO1_23_Y));
    AND2 AND2_33 (.A(\MEM_WADDR[12] ), .B(GND), .Y(AND2_33_Y));
    XOR2 XOR2_44 (.A(\WBINSYNCSHIFT[6] ), .B(INV_5_Y), .Y(XOR2_44_Y));
    DFN1C0 \DFN1C0_RGRYSYNC[2]  (.D(DFN1C0_6_Q), .CLK(WCLOCK), .CLR(
        WRITE_RESET_P), .Q(\RGRYSYNC[2] ));
    DFN1C0 \DFN1C0_RDCNT[11]  (.D(\RDIFF[11] ), .CLK(RCLOCK), .CLR(
        READ_RESET_P), .Q(RDCNT[11]));
    AO1 AO1_10 (.A(XOR2_49_Y), .B(AND2_92_Y), .C(AND2_51_Y), .Y(
        AO1_10_Y));
    XNOR3 XNOR3_49 (.A(\RGRYSYNC[3] ), .B(\RGRYSYNC[2] ), .C(XOR3_7_Y), 
        .Y(XNOR3_49_Y));
    XNOR3 XNOR3_30 (.A(\RGRYSYNC[12] ), .B(\RGRYSYNC[11] ), .C(
        \RGRYSYNC[10] ), .Y(XNOR3_30_Y));
    XOR2 XOR2_41 (.A(\WBINSYNCSHIFT[7] ), .B(INV_7_Y), .Y(XOR2_41_Y));
    XOR2 XOR2_35 (.A(\WBINNXTSHIFT[1] ), .B(\WBINNXTSHIFT[2] ), .Y(
        XOR2_35_Y));
    XNOR2 XNOR2_24 (.A(\RBINNXTSHIFT[4] ), .B(\WBINSYNCSHIFT[4] ), .Y(
        XNOR2_24_Y));
    DFN1C0 \DFN1C0_RGRYSYNC[0]  (.D(DFN1C0_27_Q), .CLK(WCLOCK), .CLR(
        WRITE_RESET_P), .Q(\RGRYSYNC[0] ));
    XOR2 \XOR2_RBINNXTSHIFT[10]  (.A(XOR2_39_Y), .B(AO1_26_Y), .Y(
        \RBINNXTSHIFT[10] ));
    XOR2 XOR2_80 (.A(\MEM_WADDR[9] ), .B(GND), .Y(XOR2_80_Y));
    DFN1C0 \DFN1C0_WGRY[1]  (.D(XOR2_35_Y), .CLK(WCLOCK), .CLR(
        WRITE_RESET_P), .Q(\WGRY[1] ));
    DFN1P0 DFN1P0_EMPTY (.D(EMPTYINT), .CLK(RCLOCK), .PRE(READ_RESET_P)
        , .Q(EMPTY));
    DFN1C0 \DFN1C0_WGRYSYNC[4]  (.D(DFN1C0_5_Q), .CLK(RCLOCK), .CLR(
        READ_RESET_P), .Q(\WGRYSYNC[4] ));
    XNOR3 XNOR3_29 (.A(\WGRYSYNC[9] ), .B(\WGRYSYNC[8] ), .C(
        \WGRYSYNC[7] ), .Y(XNOR3_29_Y));
    XNOR3 \XNOR3_RBINSYNCSHIFT[4]  (.A(XNOR3_30_Y), .B(XNOR3_41_Y), .C(
        XNOR3_9_Y), .Y(\RBINSYNCSHIFT[4] ));
    DFN1C0 DFN1C0_27 (.D(\RGRY[0] ), .CLK(WCLOCK), .CLR(WRITE_RESET_P), 
        .Q(DFN1C0_27_Q));
    XOR2 XOR2_78 (.A(\MEM_WADDR[6] ), .B(GND), .Y(XOR2_78_Y));
    XOR2 \XOR2_RDIFF[11]  (.A(XOR2_12_Y), .B(AO1_41_Y), .Y(\RDIFF[11] )
        );
    AO1 AO1_30 (.A(XOR2_81_Y), .B(AO1_36_Y), .C(AND2_71_Y), .Y(
        AO1_30_Y));
    XOR2 \XOR2_WBINSYNCSHIFT[11]  (.A(\WGRYSYNC[12] ), .B(
        \WGRYSYNC[11] ), .Y(\WBINSYNCSHIFT[11] ));
    XOR2 \XOR2_RBINNXTSHIFT[7]  (.A(XOR2_83_Y), .B(AO1_32_Y), .Y(
        \RBINNXTSHIFT[7] ));
    AND2 AND2_41 (.A(AND2_82_Y), .B(AND2_81_Y), .Y(AND2_41_Y));
    AND2 AND2_0 (.A(AND2_87_Y), .B(AND2_4_Y), .Y(AND2_0_Y));
    DFN1C0 \DFN1C0_RGRY[12]  (.D(XOR2_45_Y), .CLK(RCLOCK), .CLR(
        READ_RESET_P), .Q(\RGRY[12] ));
    XOR2 XOR2_69 (.A(\MEM_RADDR[3] ), .B(GND), .Y(XOR2_69_Y));
    AO1 AO1_16 (.A(XOR2_31_Y), .B(AND2_5_Y), .C(AND2_19_Y), .Y(
        AO1_16_Y));
    AND2 AND2_17 (.A(XOR2_79_Y), .B(XOR2_30_Y), .Y(AND2_17_Y));
    XNOR2 \XNOR2_WBINSYNCSHIFT[1]  (.A(XNOR3_28_Y), .B(XNOR3_40_Y), .Y(
        \WBINSYNCSHIFT[1] ));
    NOR2A NOR2A_0 (.A(\RBINNXTSHIFT[0] ), .B(\WBINSYNCSHIFT[0] ), .Y(
        NOR2A_0_Y));
    AO1 AO1_29 (.A(AND2_4_Y), .B(AO1_12_Y), .C(AO1_48_Y), .Y(AO1_29_Y));
    XOR2 XOR2_6 (.A(\RBINNXTSHIFT[11] ), .B(\RBINNXTSHIFT[12] ), .Y(
        XOR2_6_Y));
    AND2 AND2_77 (.A(AND2_96_Y), .B(XOR2_19_Y), .Y(AND2_77_Y));
    DFN1C0 \DFN1C0_WGRY[12]  (.D(XOR2_70_Y), .CLK(WCLOCK), .CLR(
        WRITE_RESET_P), .Q(\WGRY[12] ));
    AND2 AND2_54 (.A(AND2_41_Y), .B(XOR2_81_Y), .Y(AND2_54_Y));
    AO1 AO1_13 (.A(XOR2_94_Y), .B(AND2_74_Y), .C(AND2_50_Y), .Y(
        AO1_13_Y));
    XOR2 XOR2_93 (.A(\WBINSYNCSHIFT[6] ), .B(INV_5_Y), .Y(XOR2_93_Y));
    DFN1C0 \DFN1C0_RDCNT[10]  (.D(\RDIFF[10] ), .CLK(RCLOCK), .CLR(
        READ_RESET_P), .Q(RDCNT[10]));
    XOR2 XOR2_84 (.A(\RBINNXTSHIFT[4] ), .B(\RBINNXTSHIFT[5] ), .Y(
        XOR2_84_Y));
    XNOR3 \XNOR3_RBINSYNCSHIFT[2]  (.A(XNOR3_3_Y), .B(XNOR3_44_Y), .C(
        XNOR3_49_Y), .Y(\RBINSYNCSHIFT[2] ));
    DFN1C0 \DFN1C0_MEM_WADDR[6]  (.D(\WBINNXTSHIFT[6] ), .CLK(WCLOCK), 
        .CLR(WRITE_RESET_P), .Q(\MEM_WADDR[6] ));
    XOR2 \XOR2_WBINNXTSHIFT[5]  (.A(XOR2_53_Y), .B(AO1_30_Y), .Y(
        \WBINNXTSHIFT[5] ));
    XOR2 XOR2_81 (.A(\MEM_WADDR[4] ), .B(GND), .Y(XOR2_81_Y));
    XOR2 \XOR2_RDIFF[6]  (.A(XOR2_93_Y), .B(AO1_52_Y), .Y(\RDIFF[6] ));
    XOR2 XOR2_53 (.A(\MEM_WADDR[5] ), .B(GND), .Y(XOR2_53_Y));
    AO1 AO1_36 (.A(AND2_81_Y), .B(AO1_1_Y), .C(AO1_31_Y), .Y(AO1_36_Y));
    XNOR2 XNOR2_23 (.A(\RBINNXTSHIFT[10] ), .B(\WBINSYNCSHIFT[10] ), 
        .Y(XNOR2_23_Y));
    AND2 AND2_81 (.A(XOR2_22_Y), .B(XOR2_86_Y), .Y(AND2_81_Y));
    XOR2 \XOR2_WBINNXTSHIFT[10]  (.A(XOR2_36_Y), .B(AO1_21_Y), .Y(
        \WBINNXTSHIFT[10] ));
    DFN1C0 DFN1C0_19 (.D(\RGRY[12] ), .CLK(WCLOCK), .CLR(WRITE_RESET_P)
        , .Q(DFN1C0_19_Q));
    DFN1C0 \DFN1C0_RDCNT[4]  (.D(\RDIFF[4] ), .CLK(RCLOCK), .CLR(
        READ_RESET_P), .Q(RDCNT[4]));
    AO1 AO1_33 (.A(XOR2_34_Y), .B(AO1_22_Y), .C(AND2_33_Y), .Y(
        AO1_33_Y));
    AO1 AO1_44 (.A(XOR2_91_Y), .B(AND2_60_Y), .C(AND2_59_Y), .Y(
        AO1_44_Y));
    DFN1C0 \DFN1C0_WGRYSYNC[3]  (.D(DFN1C0_26_Q), .CLK(RCLOCK), .CLR(
        READ_RESET_P), .Q(\WGRYSYNC[3] ));
    XNOR2 XNOR2_12 (.A(\RBINNXTSHIFT[0] ), .B(\WBINSYNCSHIFT[0] ), .Y(
        XNOR2_12_Y));
    XNOR2 XNOR2_7 (.A(\RBINNXTSHIFT[1] ), .B(\WBINSYNCSHIFT[1] ), .Y(
        XNOR2_7_Y));
    XOR2 XOR2_12 (.A(\WBINSYNCSHIFT[11] ), .B(INV_8_Y), .Y(XOR2_12_Y));
    AND2 AND2_48 (.A(READDOMAIN_WMSB), .B(INV_6_Y), .Y(AND2_48_Y));
    AND2 AND2_45 (.A(\MEM_RADDR[11] ), .B(GND), .Y(AND2_45_Y));
    DFN1C0 DFN1C0_5 (.D(\WGRY[4] ), .CLK(RCLOCK), .CLR(READ_RESET_P), 
        .Q(DFN1C0_5_Q));
    DFN1C0 DFN1C0_21 (.D(\RGRY[6] ), .CLK(WCLOCK), .CLR(WRITE_RESET_P), 
        .Q(DFN1C0_21_Q));
    AO1 AO1_19 (.A(AND2_30_Y), .B(AO1_23_Y), .C(AO1_13_Y), .Y(AO1_19_Y)
        );
    XOR2 \XOR2_WBINNXTSHIFT[7]  (.A(XOR2_33_Y), .B(AO1_18_Y), .Y(
        \WBINNXTSHIFT[7] ));
    DFN1C0 \DFN1C0_MEM_RADDR[12]  (.D(\RBINNXTSHIFT[12] ), .CLK(RCLOCK)
        , .CLR(READ_RESET_P), .Q(\MEM_RADDR[12] ));
    XOR2 XOR2_26 (.A(\WBINSYNCSHIFT[11] ), .B(INV_8_Y), .Y(XOR2_26_Y));
    DFN1C0 DFN1C0_1 (.D(\RGRY[9] ), .CLK(WCLOCK), .CLR(WRITE_RESET_P), 
        .Q(DFN1C0_1_Q));
    AND2 AND2_59 (.A(\WBINSYNCSHIFT[10] ), .B(INV_11_Y), .Y(AND2_59_Y));
    DFN1C0 \DFN1C0_RGRY[10]  (.D(XOR2_87_Y), .CLK(RCLOCK), .CLR(
        READ_RESET_P), .Q(\RGRY[10] ));
    XOR2 \XOR2_RDIFF[4]  (.A(XOR2_64_Y), .B(AO1_53_Y), .Y(\RDIFF[4] ));
    DFN1C0 \DFN1C0_WGRYSYNC[7]  (.D(DFN1C0_8_Q), .CLK(RCLOCK), .CLR(
        READ_RESET_P), .Q(\WGRYSYNC[7] ));
    AND2 AND2_4 (.A(AND2_27_Y), .B(AND2_44_Y), .Y(AND2_4_Y));
    XOR2 XOR2_90 (.A(\MEM_WADDR[3] ), .B(GND), .Y(XOR2_90_Y));
    AND2 AND2_FULLINT (.A(AND3_1_Y), .B(XOR2_55_Y), .Y(FULLINT));
    DFN1C0 \DFN1C0_RDCNT[3]  (.D(\RDIFF[3] ), .CLK(RCLOCK), .CLR(
        READ_RESET_P), .Q(RDCNT[3]));
    AO1 AO1_39 (.A(XOR2_25_Y), .B(AO1_9_Y), .C(AND2_85_Y), .Y(AO1_39_Y)
        );
    AND2 AND2_40 (.A(AND2_52_Y), .B(XOR2_71_Y), .Y(AND2_40_Y));
    XNOR3 XNOR3_12 (.A(\RGRYSYNC[3] ), .B(\RGRYSYNC[2] ), .C(
        \RGRYSYNC[1] ), .Y(XNOR3_12_Y));
    AND2 AND2_88 (.A(XOR2_14_Y), .B(XOR2_91_Y), .Y(AND2_88_Y));
    AND2 AND2_85 (.A(\MEM_WADDR[8] ), .B(GND), .Y(AND2_85_Y));
    XOR2 XOR2_50 (.A(\MEM_RADDR[1] ), .B(GND), .Y(XOR2_50_Y));
    DFN1C0 \DFN1C0_WGRYSYNC[6]  (.D(DFN1C0_20_Q), .CLK(RCLOCK), .CLR(
        READ_RESET_P), .Q(\WGRYSYNC[6] ));
    AND2 AND2_94 (.A(AND2_0_Y), .B(AND2_83_Y), .Y(AND2_94_Y));
    AND2 AND2_42 (.A(XOR2_26_Y), .B(XOR2_82_Y), .Y(AND2_42_Y));
    DFN1C0 \DFN1C0_WGRY[8]  (.D(XOR2_62_Y), .CLK(WCLOCK), .CLR(
        WRITE_RESET_P), .Q(\WGRY[8] ));
    XNOR2 XNOR2_5 (.A(\RBINSYNCSHIFT[5] ), .B(\WBINNXTSHIFT[5] ), .Y(
        XNOR2_5_Y));
    AO1 AO1_5 (.A(AND2_80_Y), .B(AO1_2_Y), .C(AO1_19_Y), .Y(AO1_5_Y));
    AND2 AND2_67 (.A(INV_0_Y), .B(INV_4_Y), .Y(AND2_67_Y));
    XNOR2 XNOR2_16 (.A(\RBINNXTSHIFT[8] ), .B(\WBINSYNCSHIFT[8] ), .Y(
        XNOR2_16_Y));
    XOR2 \XOR2_RBINSYNCSHIFT[11]  (.A(\RGRYSYNC[12] ), .B(
        \RGRYSYNC[11] ), .Y(\RBINSYNCSHIFT[11] ));
    XNOR3 XNOR3_41 (.A(\RGRYSYNC[9] ), .B(\RGRYSYNC[8] ), .C(
        \RGRYSYNC[7] ), .Y(XNOR3_41_Y));
    XNOR3 XNOR3_32 (.A(\WGRYSYNC[6] ), .B(\WGRYSYNC[5] ), .C(
        \WGRYSYNC[4] ), .Y(XNOR3_32_Y));
    DFN1C0 \DFN1C0_RGRY[3]  (.D(XOR2_58_Y), .CLK(RCLOCK), .CLR(
        READ_RESET_P), .Q(\RGRY[3] ));
    XOR2 XOR2_94 (.A(\WBINSYNCSHIFT[8] ), .B(INV_1_Y), .Y(XOR2_94_Y));
    XOR3 XOR3_2 (.A(\RGRYSYNC[12] ), .B(\RGRYSYNC[11] ), .C(
        \RGRYSYNC[10] ), .Y(XOR3_2_Y));
    XOR2 XOR2_39 (.A(\MEM_RADDR[10] ), .B(GND), .Y(XOR2_39_Y));
    AND2 AND2_8 (.A(XOR2_19_Y), .B(XOR2_44_Y), .Y(AND2_8_Y));
    XOR2 XOR2_91 (.A(\WBINSYNCSHIFT[10] ), .B(INV_11_Y), .Y(XOR2_91_Y));
    AND2 AND2_80 (.A(AND2_8_Y), .B(AND2_30_Y), .Y(AND2_80_Y));
    XNOR2 \XNOR2_WBINSYNCSHIFT[9]  (.A(\WGRYSYNC[9] ), .B(XNOR3_22_Y), 
        .Y(\WBINSYNCSHIFT[9] ));
    XOR2 XOR2_3 (.A(\WBINNXTSHIFT[11] ), .B(\WBINNXTSHIFT[12] ), .Y(
        XOR2_3_Y));
    XOR2 XOR2_54 (.A(\WBINNXTSHIFT[10] ), .B(\WBINNXTSHIFT[11] ), .Y(
        XOR2_54_Y));
    XNOR3 XNOR3_21 (.A(\WGRYSYNC[12] ), .B(\WGRYSYNC[11] ), .C(
        \WGRYSYNC[10] ), .Y(XNOR3_21_Y));
    XOR3 XOR3_1 (.A(\RGRYSYNC[12] ), .B(\RGRYSYNC[11] ), .C(
        \RGRYSYNC[10] ), .Y(XOR3_1_Y));
    XOR2 \XOR2_RBINNXTSHIFT[11]  (.A(XOR2_100_Y), .B(AO1_54_Y), .Y(
        \RBINNXTSHIFT[11] ));
    XOR2 XOR2_51 (.A(\WBINSYNCSHIFT[3] ), .B(INV_2_Y), .Y(XOR2_51_Y));
    AO1 AO1_27 (.A(XOR2_56_Y), .B(AND2_85_Y), .C(AND2_73_Y), .Y(
        AO1_27_Y));
    AND2 AND2_82 (.A(XOR2_47_Y), .B(XOR2_40_Y), .Y(AND2_82_Y));
    XOR2 XOR2_66 (.A(\MEM_WADDR[1] ), .B(GND), .Y(XOR2_66_Y));
    DFN1C0 DFN1C0_24 (.D(\WGRY[5] ), .CLK(RCLOCK), .CLR(READ_RESET_P), 
        .Q(DFN1C0_24_Q));
    AND2 AND2_56 (.A(AND2_0_Y), .B(XOR2_20_Y), .Y(AND2_56_Y));
    XNOR3 \XNOR3_RBINSYNCSHIFT[0]  (.A(XNOR3_43_Y), .B(XNOR3_12_Y), .C(
        XNOR3_5_Y), .Y(\RBINSYNCSHIFT[0] ));
    INV INV_10 (.A(\RBINNXTSHIFT[5] ), .Y(INV_10_Y));
    DFN1C0 \DFN1C0_MEM_WADDR[1]  (.D(\WBINNXTSHIFT[1] ), .CLK(WCLOCK), 
        .CLR(WRITE_RESET_P), .Q(\MEM_WADDR[1] ));
    XNOR3 XNOR3_16 (.A(\WGRYSYNC[6] ), .B(\WGRYSYNC[5] ), .C(
        \WGRYSYNC[4] ), .Y(XNOR3_16_Y));
    XOR2 \XOR2_RBINNXTSHIFT[1]  (.A(XOR2_50_Y), .B(AND2_91_Y), .Y(
        \RBINNXTSHIFT[1] ));
    DFN1C0 \DFN1C0_RDCNT[9]  (.D(\RDIFF[9] ), .CLK(RCLOCK), .CLR(
        READ_RESET_P), .Q(RDCNT[9]));
    XOR2 XOR2_17 (.A(\MEM_WADDR[12] ), .B(GND), .Y(XOR2_17_Y));
    XOR2 XOR2_73 (.A(\WBINNXTSHIFT[3] ), .B(\WBINNXTSHIFT[4] ), .Y(
        XOR2_73_Y));
    AND2 AND2_53 (.A(\WBINSYNCSHIFT[5] ), .B(INV_10_Y), .Y(AND2_53_Y));
    DFN1C0 DFN1C0_13 (.D(\WGRY[0] ), .CLK(RCLOCK), .CLR(READ_RESET_P), 
        .Q(DFN1C0_13_Q));
    XNOR3 XNOR3_51 (.A(\RGRYSYNC[9] ), .B(\RGRYSYNC[8] ), .C(
        \RGRYSYNC[7] ), .Y(XNOR3_51_Y));
    AND3 AND3_7 (.A(XNOR2_12_Y), .B(XNOR2_7_Y), .C(XNOR2_13_Y), .Y(
        AND3_7_Y));
    XOR2 XOR2_28 (.A(\RBINNXTSHIFT[1] ), .B(\RBINNXTSHIFT[2] ), .Y(
        XOR2_28_Y));
    INV INV_9 (.A(\RBINNXTSHIFT[2] ), .Y(INV_9_Y));
    XNOR3 XNOR3_36 (.A(XNOR3_37_Y), .B(XNOR3_7_Y), .C(XNOR3_19_Y), .Y(
        XNOR3_36_Y));
    DFN1C0 \DFN1C0_MEM_WADDR[5]  (.D(\WBINNXTSHIFT[5] ), .CLK(WCLOCK), 
        .CLR(WRITE_RESET_P), .Q(\MEM_WADDR[5] ));
    XOR2 XOR2_15 (.A(\MEM_RADDR[4] ), .B(GND), .Y(XOR2_15_Y));
    XNOR3 XNOR3_48 (.A(\WGRYSYNC[9] ), .B(\WGRYSYNC[8] ), .C(
        \WGRYSYNC[7] ), .Y(XNOR3_48_Y));
    XOR2 \XOR2_RDIFF[5]  (.A(XOR2_29_Y), .B(AO1_2_Y), .Y(\RDIFF[5] ));
    DFN1C0 \DFN1C0_MEM_RADDR[0]  (.D(\RBINNXTSHIFT[0] ), .CLK(RCLOCK), 
        .CLR(READ_RESET_P), .Q(\MEM_RADDR[0] ));
    AO1 AO1_17 (.A(AND2_86_Y), .B(AO1_36_Y), .C(AO1_7_Y), .Y(AO1_17_Y));
    XNOR3 \XNOR3_WBINSYNCSHIFT[4]  (.A(XNOR3_4_Y), .B(XNOR3_13_Y), .C(
        XNOR3_32_Y), .Y(\WBINSYNCSHIFT[4] ));
    XNOR2 XNOR2_17 (.A(\RBINSYNCSHIFT[1] ), .B(\WBINNXTSHIFT[1] ), .Y(
        XNOR2_17_Y));
    DFN1C0 \DFN1C0_MEM_RADDR[10]  (.D(\RBINNXTSHIFT[10] ), .CLK(RCLOCK)
        , .CLR(READ_RESET_P), .Q(\MEM_RADDR[10] ));
    XOR2 \XOR2_WBINNXTSHIFT[11]  (.A(XOR2_67_Y), .B(AO1_42_Y), .Y(
        \WBINNXTSHIFT[11] ));
    AND3 AND3_4 (.A(XNOR2_15_Y), .B(XNOR2_8_Y), .C(XNOR2_2_Y), .Y(
        AND3_4_Y));
    XNOR3 XNOR3_28 (.A(\WGRYSYNC[3] ), .B(\WGRYSYNC[2] ), .C(
        \WGRYSYNC[1] ), .Y(XNOR3_28_Y));
    DFN1C0 \DFN1C0_RGRY[0]  (.D(XOR2_18_Y), .CLK(RCLOCK), .CLR(
        READ_RESET_P), .Q(\RGRY[0] ));
    XOR2 \XOR2_WBINNXTSHIFT[1]  (.A(XOR2_66_Y), .B(AND2_39_Y), .Y(
        \WBINNXTSHIFT[1] ));
    AND2 AND2_21 (.A(XOR2_0_Y), .B(XOR2_49_Y), .Y(AND2_21_Y));
    XOR3 XOR3_7 (.A(\RGRYSYNC[12] ), .B(\RGRYSYNC[11] ), .C(
        \RGRYSYNC[10] ), .Y(XOR3_7_Y));
    AO1 AO1_37 (.A(XOR2_22_Y), .B(AO1_1_Y), .C(AND2_13_Y), .Y(AO1_37_Y)
        );
    DFN1C0 \DFN1C0_WGRY[4]  (.D(XOR2_63_Y), .CLK(WCLOCK), .CLR(
        WRITE_RESET_P), .Q(\WGRY[4] ));
    DFN1C0 DFN1C0_25 (.D(\RGRY[8] ), .CLK(WCLOCK), .CLR(WRITE_RESET_P), 
        .Q(DFN1C0_25_Q));
    XNOR3 XNOR3_17 (.A(\WGRYSYNC[12] ), .B(\WGRYSYNC[11] ), .C(
        \WGRYSYNC[10] ), .Y(XNOR3_17_Y));
    XOR2 XOR2_0 (.A(\WBINSYNCSHIFT[3] ), .B(INV_2_Y), .Y(XOR2_0_Y));
    NAND2 NAND2_1 (.A(EMPTY), .B(VCC), .Y(NAND2_1_Y));
    XOR2 XOR2_70 (.A(\WBINNXTSHIFT[12] ), .B(GND), .Y(XOR2_70_Y));
    AND2 AND2_96 (.A(AND2_12_Y), .B(AND2_21_Y), .Y(AND2_96_Y));
    DFN1C0 DFN1C0_22 (.D(\WGRY[9] ), .CLK(RCLOCK), .CLR(READ_RESET_P), 
        .Q(DFN1C0_22_Q));
    XNOR3 \XNOR3_WBINSYNCSHIFT[6]  (.A(\WGRYSYNC[6] ), .B(XOR3_3_Y), 
        .C(XNOR3_26_Y), .Y(\WBINSYNCSHIFT[6] ));
    DFN1C0 \DFN1C0_RGRYSYNC[8]  (.D(DFN1C0_25_Q), .CLK(WCLOCK), .CLR(
        WRITE_RESET_P), .Q(\RGRYSYNC[8] ));
    AO1 AO1_4 (.A(XOR2_11_Y), .B(OR3_0_Y), .C(AND2_55_Y), .Y(AO1_4_Y));
    XOR2 XOR2_68 (.A(\MEM_RADDR[10] ), .B(GND), .Y(XOR2_68_Y));
    AND2 AND2_37 (.A(\WBINSYNCSHIFT[1] ), .B(INV_0_Y), .Y(AND2_37_Y));
    XNOR3 XNOR3_4 (.A(\WGRYSYNC[12] ), .B(\WGRYSYNC[11] ), .C(
        \WGRYSYNC[10] ), .Y(XNOR3_4_Y));
    AND2 AND2_93 (.A(AND2_95_Y), .B(XOR2_68_Y), .Y(AND2_93_Y));
    XNOR2 XNOR2_14 (.A(\RBINNXTSHIFT[3] ), .B(\WBINSYNCSHIFT[3] ), .Y(
        XNOR2_14_Y));
    XOR2 \XOR2_RBINNXTSHIFT[2]  (.A(XOR2_46_Y), .B(AO1_24_Y), .Y(
        \RBINNXTSHIFT[2] ));
    XOR2 XOR2_42 (.A(\WBINNXTSHIFT[0] ), .B(\WBINNXTSHIFT[1] ), .Y(
        XOR2_42_Y));
    XNOR3 XNOR3_37 (.A(\RGRYSYNC[12] ), .B(\RGRYSYNC[11] ), .C(
        \RGRYSYNC[10] ), .Y(XNOR3_37_Y));
    AO1 AO1_21 (.A(AND2_11_Y), .B(AO1_9_Y), .C(AO1_27_Y), .Y(AO1_21_Y));
    DFN1C0 \DFN1C0_MEM_RADDR[9]  (.D(\RBINNXTSHIFT[9] ), .CLK(RCLOCK), 
        .CLR(READ_RESET_P), .Q(\MEM_RADDR[9] ));
    XOR2 XOR2_36 (.A(\MEM_WADDR[10] ), .B(GND), .Y(XOR2_36_Y));
    XOR2 XOR2_74 (.A(\RBINNXTSHIFT[8] ), .B(\RBINNXTSHIFT[9] ), .Y(
        XOR2_74_Y));
    XNOR3 \XNOR3_RBINSYNCSHIFT[6]  (.A(\RGRYSYNC[6] ), .B(XOR3_5_Y), 
        .C(XNOR3_0_Y), .Y(\RBINSYNCSHIFT[6] ));
    XNOR2 XNOR2_8 (.A(\RBINSYNCSHIFT[7] ), .B(\WBINNXTSHIFT[7] ), .Y(
        XNOR2_8_Y));
    XNOR3 XNOR3_2 (.A(\RGRYSYNC[3] ), .B(\RGRYSYNC[2] ), .C(
        \RGRYSYNC[1] ), .Y(XNOR3_2_Y));
    XOR2 XOR2_71 (.A(\MEM_RADDR[6] ), .B(GND), .Y(XOR2_71_Y));
    AND2 AND2_28 (.A(AND2_41_Y), .B(AND2_86_Y), .Y(AND2_28_Y));
    AND2 AND2_25 (.A(XNOR2_23_Y), .B(XNOR2_4_Y), .Y(AND2_25_Y));
    AO1 AO1_48 (.A(AND2_44_Y), .B(AO1_16_Y), .C(AO1_55_Y), .Y(AO1_48_Y)
        );
    DFN1C0 \DFN1C0_RDCNT[6]  (.D(\RDIFF[6] ), .CLK(RCLOCK), .CLR(
        READ_RESET_P), .Q(RDCNT[6]));
    DFN1C0 \DFN1C0_MEM_RADDR[11]  (.D(\RBINNXTSHIFT[11] ), .CLK(RCLOCK)
        , .CLR(READ_RESET_P), .Q(\MEM_RADDR[11] ));
    DFN1C0 \DFN1C0_WGRYSYNC[5]  (.D(DFN1C0_24_Q), .CLK(RCLOCK), .CLR(
        READ_RESET_P), .Q(\WGRYSYNC[5] ));
    GND GND_power_inst1 (.Y(GND_power_net1));
    VCC VCC_power_inst1 (.Y(VCC_power_net1));
    
endmodule

// _Disclaimer: Please leave the following comments in the file, they are for internal purposes only._


// _GEN_File_Contents_

// Version:11.9.5.5
// ACTGENU_CALL:1
// BATCH:T
// FAM:PA3LCLP
// OUTFORMAT:Verilog
// LPMTYPE:LPM_SOFTFIFO
// LPM_HINT:MEMFF
// INSERT_PAD:NO
// INSERT_IOREG:NO
// GEN_BHV_VHDL_VAL:F
// GEN_BHV_VERILOG_VAL:F
// MGNTIMER:F
// MGNCMPL:T
// DESDIR:C:/Microsemi/earEEG_prototype_vivado/smartgen\fifo_1b_1b
// GEN_BEHV_MODULE:F
// SMARTGEN_DIE:IS6X6M2LP
// SMARTGEN_PACKAGE:fg144
// AGENIII_IS_SUBPROJECT_LIBERO:T
// WWIDTH:1
// WDEPTH:4096
// RWIDTH:1
// RDEPTH:4096
// CLKS:2
// WCLOCK_PN:WCLOCK
// RCLOCK_PN:RCLOCK
// WCLK_EDGE:RISE
// RCLK_EDGE:RISE
// ACLR_PN:RESET
// RESET_POLARITY:1
// INIT_RAM:F
// WE_POLARITY:1
// RE_POLARITY:1
// FF_PN:FULL
// AF_PN:AFULL
// WACK_PN:WACK
// OVRFLOW_PN:OVERFLOW
// WRCNT_PN:WRCNT
// WE_PN:WE
// EF_PN:EMPTY
// AE_PN:AEMPTY
// DVLD_PN:DVLD
// UDRFLOW_PN:UNDERFLOW
// RDCNT_PN:RDCNT
// RE_PN:RE
// CONTROLLERONLY:F
// FSTOP:YES
// ESTOP:YES
// WRITEACK:NO
// OVERFLOW:NO
// WRCOUNT:NO
// DATAVALID:NO
// UNDERFLOW:NO
// RDCOUNT:YES
// AF_PORT_PN:AFVAL
// AE_PORT_PN:AEVAL
// AFFLAG:NONE
// AEFLAG:NONE
// DATA_IN_PN:DATA
// DATA_OUT_PN:Q
// CASCADE:1

// _End_Comments_

